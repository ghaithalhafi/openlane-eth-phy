VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter32
  CLASS BLOCK ;
  FOREIGN counter32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 96.520 BY 107.240 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 95.440 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 95.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END clk
  PIN count[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END count[0]
  PIN count[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END count[10]
  PIN count[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END count[11]
  PIN count[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END count[12]
  PIN count[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END count[13]
  PIN count[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END count[14]
  PIN count[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END count[15]
  PIN count[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END count[16]
  PIN count[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END count[17]
  PIN count[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END count[18]
  PIN count[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END count[19]
  PIN count[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END count[1]
  PIN count[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 103.240 45.450 107.240 ;
    END
  END count[20]
  PIN count[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 103.240 42.230 107.240 ;
    END
  END count[21]
  PIN count[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 103.240 55.110 107.240 ;
    END
  END count[22]
  PIN count[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 103.240 58.330 107.240 ;
    END
  END count[23]
  PIN count[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.520 44.240 96.520 44.840 ;
    END
  END count[24]
  PIN count[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.520 40.840 96.520 41.440 ;
    END
  END count[25]
  PIN count[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.520 47.640 96.520 48.240 ;
    END
  END count[26]
  PIN count[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.520 51.040 96.520 51.640 ;
    END
  END count[27]
  PIN count[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.520 68.040 96.520 68.640 ;
    END
  END count[28]
  PIN count[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.520 71.440 96.520 72.040 ;
    END
  END count[29]
  PIN count[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END count[2]
  PIN count[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.520 64.640 96.520 65.240 ;
    END
  END count[30]
  PIN count[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.520 61.240 96.520 61.840 ;
    END
  END count[31]
  PIN count[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END count[3]
  PIN count[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END count[4]
  PIN count[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END count[5]
  PIN count[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END count[6]
  PIN count[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END count[7]
  PIN count[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END count[8]
  PIN count[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END count[9]
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END en
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 92.520 20.440 96.520 21.040 ;
    END
  END rst_n
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 90.810 95.390 ;
      LAYER li1 ;
        RECT 5.520 10.795 90.620 95.285 ;
      LAYER met1 ;
        RECT 4.210 10.640 90.620 95.440 ;
      LAYER met2 ;
        RECT 4.230 102.960 41.670 103.770 ;
        RECT 42.510 102.960 44.890 103.770 ;
        RECT 45.730 102.960 54.550 103.770 ;
        RECT 55.390 102.960 57.770 103.770 ;
        RECT 58.610 102.960 89.150 103.770 ;
        RECT 4.230 4.280 89.150 102.960 ;
        RECT 4.230 4.000 15.910 4.280 ;
        RECT 16.750 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.210 4.280 ;
        RECT 65.050 4.000 89.150 4.280 ;
      LAYER met3 ;
        RECT 3.990 72.440 92.520 95.365 ;
        RECT 4.400 71.040 92.120 72.440 ;
        RECT 3.990 69.040 92.520 71.040 ;
        RECT 4.400 67.640 92.120 69.040 ;
        RECT 3.990 65.640 92.520 67.640 ;
        RECT 4.400 64.240 92.120 65.640 ;
        RECT 3.990 62.240 92.520 64.240 ;
        RECT 4.400 60.840 92.120 62.240 ;
        RECT 3.990 58.840 92.520 60.840 ;
        RECT 4.400 57.440 92.520 58.840 ;
        RECT 3.990 52.040 92.520 57.440 ;
        RECT 4.400 50.640 92.120 52.040 ;
        RECT 3.990 48.640 92.520 50.640 ;
        RECT 3.990 47.240 92.120 48.640 ;
        RECT 3.990 45.240 92.520 47.240 ;
        RECT 3.990 43.840 92.120 45.240 ;
        RECT 3.990 41.840 92.520 43.840 ;
        RECT 4.400 40.440 92.120 41.840 ;
        RECT 3.990 38.440 92.520 40.440 ;
        RECT 4.400 37.040 92.520 38.440 ;
        RECT 3.990 35.040 92.520 37.040 ;
        RECT 4.400 33.640 92.520 35.040 ;
        RECT 3.990 21.440 92.520 33.640 ;
        RECT 3.990 20.040 92.120 21.440 ;
        RECT 3.990 6.295 92.520 20.040 ;
      LAYER met4 ;
        RECT 41.695 6.295 42.025 41.985 ;
  END
END counter32
END LIBRARY

