* NGSPICE file created from eth_phy_1g.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

.subckt eth_phy_1g VGND VPWR clk eth_data_in[0] eth_data_in[1] eth_data_in[2] eth_data_in[3]
+ eth_data_in[4] eth_data_in[5] eth_data_in[6] eth_data_in[7] eth_valid_in phy_data_out[0]
+ phy_data_out[1] phy_data_out[2] phy_data_out[3] phy_data_out[4] phy_data_out[5]
+ phy_data_out[6] phy_data_out[7] phy_data_out[8] phy_data_out[9] phy_valid_out rst
X_49_ net10 VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__inv_2
Xoutput20 net20 VGND VGND VPWR VPWR phy_data_out[9] sky130_fd_sc_hd__buf_2
X_65_ net20 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_4_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_48_ net10 VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__inv_2
Xoutput21 net21 VGND VGND VPWR VPWR phy_valid_out sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_64_ net20 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_47_ net10 VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__inv_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput11 net11 VGND VGND VPWR VPWR phy_data_out[0] sky130_fd_sc_hd__buf_2
X_63_ net19 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_46_ _22_ _26_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_5_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput12 net12 VGND VGND VPWR VPWR phy_data_out[1] sky130_fd_sc_hd__buf_2
X_29_ net28 VGND VGND VPWR VPWR _17_ sky130_fd_sc_hd__inv_2
X_62_ net17 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_8_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_45_ _16_ u_pcs.rd_pos VGND VGND VPWR VPWR _26_ sky130_fd_sc_hd__and2_1
X_28_ net9 VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__inv_2
Xoutput13 net13 VGND VGND VPWR VPWR phy_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_61_ clknet_1_1__leaf_clk _14_ _07_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
X_44_ _16_ net25 _19_ _25_ VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__a22o_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_27_ net27 VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__inv_2
Xoutput14 net14 VGND VGND VPWR VPWR phy_data_out[3] sky130_fd_sc_hd__buf_2
X_60_ clknet_1_1__leaf_clk _13_ _06_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_1
X_43_ _22_ _21_ net1 VGND VGND VPWR VPWR _25_ sky130_fd_sc_hd__mux2_1
Xoutput15 net15 VGND VGND VPWR VPWR phy_data_out[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_42_ _16_ net23 _20_ _24_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__a211o_1
XFILLER_4_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput16 net16 VGND VGND VPWR VPWR phy_data_out[5] sky130_fd_sc_hd__buf_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_41_ _16_ _23_ VGND VGND VPWR VPWR _24_ sky130_fd_sc_hd__nor2_1
Xoutput17 net17 VGND VGND VPWR VPWR phy_data_out[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_40_ u_pcs.rd_pos net2 VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput18 net18 VGND VGND VPWR VPWR phy_data_out[7] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput19 net19 VGND VGND VPWR VPWR phy_data_out[8] sky130_fd_sc_hd__buf_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 eth_data_in[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_7_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 eth_data_in[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
Xinput3 eth_data_in[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 eth_data_in[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
Xinput5 eth_data_in[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_59_ clknet_1_0__leaf_clk _12_ _05_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
X_58_ clknet_1_0__leaf_clk _11_ _04_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Left_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 eth_data_in[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 eth_data_in[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_57_ clknet_1_0__leaf_clk _10_ _03_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
Xinput10 net22 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_4
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 eth_data_in[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_56_ clknet_1_1__leaf_clk _09_ _02_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_39_ _16_ net24 _20_ _22_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__a211o_1
Xinput9 eth_valid_in VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_55_ clknet_1_1__leaf_clk net9 _01_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_1
X_38_ _16_ _17_ _20_ _22_ VGND VGND VPWR VPWR _12_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 rst VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
X_54_ clknet_1_0__leaf_clk _08_ _00_ VGND VGND VPWR VPWR u_pcs.rd_pos sky130_fd_sc_hd__dfrtp_1
X_37_ u_pcs.rd_pos net9 VGND VGND VPWR VPWR _22_ sky130_fd_sc_hd__and2b_1
Xhold2 net12 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_1_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_53_ net10 VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__inv_2
X_36_ _16_ net26 _20_ _21_ VGND VGND VPWR VPWR _13_ sky130_fd_sc_hd__a211o_1
Xhold3 net14 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
X_52_ net10 VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__inv_2
X_35_ _15_ _16_ _20_ _21_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__a211oi_1
Xhold4 net11 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
X_51_ net10 VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__inv_2
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_34_ net9 u_pcs.rd_pos VGND VGND VPWR VPWR _21_ sky130_fd_sc_hd__and2_1
Xhold5 net20 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
X_33_ net4 net3 _18_ net9 VGND VGND VPWR VPWR _20_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_1_Left_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_50_ net10 VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__inv_2
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 net19 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ net4 net3 _18_ VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__nor3_1
Xhold7 net17 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
X_31_ net6 net5 net8 net7 VGND VGND VPWR VPWR _18_ sky130_fd_sc_hd__or4_1
XFILLER_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_30_ net10 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_5_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

