magic
tech sky130A
magscale 1 2
timestamp 1770945975
<< checkpaint >>
rect -3932 -3932 11999 14143
<< viali >>
rect 2053 7497 2087 7531
rect 2881 7497 2915 7531
rect 3525 7497 3559 7531
rect 1777 7361 1811 7395
rect 1869 7361 1903 7395
rect 2145 7361 2179 7395
rect 2605 7361 2639 7395
rect 2697 7361 2731 7395
rect 3065 7361 3099 7395
rect 3341 7361 3375 7395
rect 3801 7361 3835 7395
rect 5825 7361 5859 7395
rect 5917 7361 5951 7395
rect 6377 7361 6411 7395
rect 2421 7225 2455 7259
rect 3249 7225 3283 7259
rect 6561 7225 6595 7259
rect 1593 7157 1627 7191
rect 2329 7157 2363 7191
rect 5089 7157 5123 7191
rect 5641 7157 5675 7191
rect 6101 7157 6135 7191
rect 1869 6953 1903 6987
rect 4537 6885 4571 6919
rect 5365 6885 5399 6919
rect 1777 6817 1811 6851
rect 4905 6817 4939 6851
rect 1685 6749 1719 6783
rect 1961 6749 1995 6783
rect 2237 6749 2271 6783
rect 2605 6749 2639 6783
rect 2881 6749 2915 6783
rect 2973 6749 3007 6783
rect 3157 6749 3191 6783
rect 3249 6749 3283 6783
rect 3617 6749 3651 6783
rect 4353 6749 4387 6783
rect 4721 6749 4755 6783
rect 4813 6749 4847 6783
rect 4997 6749 5031 6783
rect 5273 6749 5307 6783
rect 5917 6749 5951 6783
rect 2329 6681 2363 6715
rect 2421 6681 2455 6715
rect 3801 6681 3835 6715
rect 5181 6681 5215 6715
rect 5641 6681 5675 6715
rect 1501 6613 1535 6647
rect 2053 6613 2087 6647
rect 2697 6613 2731 6647
rect 3433 6613 3467 6647
rect 5549 6613 5583 6647
rect 6561 6613 6595 6647
rect 1501 6409 1535 6443
rect 3709 6409 3743 6443
rect 6469 6409 6503 6443
rect 2145 6341 2179 6375
rect 4721 6341 4755 6375
rect 1501 6273 1535 6307
rect 1593 6273 1627 6307
rect 4445 6273 4479 6307
rect 6561 6273 6595 6307
rect 1777 6205 1811 6239
rect 1869 6205 1903 6239
rect 4261 6205 4295 6239
rect 6193 6205 6227 6239
rect 3617 6069 3651 6103
rect 1501 5865 1535 5899
rect 3801 5865 3835 5899
rect 3617 5797 3651 5831
rect 1869 5729 1903 5763
rect 4445 5729 4479 5763
rect 4813 5729 4847 5763
rect 1685 5661 1719 5695
rect 2145 5593 2179 5627
rect 4169 5593 4203 5627
rect 5089 5593 5123 5627
rect 4261 5525 4295 5559
rect 6561 5525 6595 5559
rect 1501 5321 1535 5355
rect 1777 5321 1811 5355
rect 2053 5321 2087 5355
rect 2513 5321 2547 5355
rect 2789 5321 2823 5355
rect 3065 5321 3099 5355
rect 5457 5321 5491 5355
rect 1685 5185 1719 5219
rect 1961 5185 1995 5219
rect 2237 5185 2271 5219
rect 2329 5185 2363 5219
rect 2881 5185 2915 5219
rect 3157 5185 3191 5219
rect 3249 5185 3283 5219
rect 5273 5185 5307 5219
rect 6561 5185 6595 5219
rect 6193 5117 6227 5151
rect 4537 4981 4571 5015
rect 5549 4981 5583 5015
rect 6469 4981 6503 5015
rect 4261 4777 4295 4811
rect 4169 4709 4203 4743
rect 4353 4709 4387 4743
rect 5641 4709 5675 4743
rect 5917 4641 5951 4675
rect 3157 4573 3191 4607
rect 3617 4573 3651 4607
rect 3801 4573 3835 4607
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 4997 4573 5031 4607
rect 5457 4573 5491 4607
rect 6469 4573 6503 4607
rect 3341 4505 3375 4539
rect 2973 4437 3007 4471
rect 3525 4437 3559 4471
rect 5181 4437 5215 4471
rect 3433 4233 3467 4267
rect 3893 4165 3927 4199
rect 2697 4097 2731 4131
rect 2973 4097 3007 4131
rect 3065 4097 3099 4131
rect 3249 4097 3283 4131
rect 3341 4097 3375 4131
rect 3617 4097 3651 4131
rect 4077 4097 4111 4131
rect 4261 4097 4295 4131
rect 6377 4097 6411 4131
rect 6469 4097 6503 4131
rect 2053 4029 2087 4063
rect 3801 4029 3835 4063
rect 4445 4029 4479 4063
rect 4721 4029 4755 4063
rect 4169 3961 4203 3995
rect 4353 3961 4387 3995
rect 2789 3893 2823 3927
rect 6193 3893 6227 3927
rect 3617 3689 3651 3723
rect 6377 3689 6411 3723
rect 1501 3621 1535 3655
rect 1869 3553 1903 3587
rect 4353 3553 4387 3587
rect 1685 3485 1719 3519
rect 3801 3485 3835 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 6561 3485 6595 3519
rect 2145 3417 2179 3451
rect 4629 3417 4663 3451
rect 3893 3349 3927 3383
rect 4169 3349 4203 3383
rect 6101 3349 6135 3383
rect 1593 3145 1627 3179
rect 3525 3145 3559 3179
rect 4905 3145 4939 3179
rect 6469 3145 6503 3179
rect 3065 3077 3099 3111
rect 3617 3009 3651 3043
rect 4077 3009 4111 3043
rect 4353 3009 4387 3043
rect 4445 3009 4479 3043
rect 4629 3009 4663 3043
rect 4721 3009 4755 3043
rect 5365 3009 5399 3043
rect 6101 3009 6135 3043
rect 6377 3009 6411 3043
rect 3341 2941 3375 2975
rect 3709 2941 3743 2975
rect 3985 2941 4019 2975
rect 5457 2941 5491 2975
rect 5181 2805 5215 2839
rect 3249 2601 3283 2635
rect 5089 2601 5123 2635
rect 5641 2601 5675 2635
rect 6101 2601 6135 2635
rect 6469 2601 6503 2635
rect 3617 2533 3651 2567
rect 3341 2397 3375 2431
rect 3433 2397 3467 2431
rect 3801 2397 3835 2431
rect 5825 2397 5859 2431
rect 5917 2397 5951 2431
rect 6377 2397 6411 2431
<< metal1 >>
rect 1104 7642 6900 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 6900 7642
rect 1104 7568 6900 7590
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7497 2099 7531
rect 2041 7491 2099 7497
rect 1946 7460 1952 7472
rect 1780 7432 1952 7460
rect 1780 7401 1808 7432
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 2056 7460 2084 7491
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 2869 7531 2927 7537
rect 2869 7528 2881 7531
rect 2648 7500 2881 7528
rect 2648 7488 2654 7500
rect 2869 7497 2881 7500
rect 2915 7497 2927 7531
rect 2869 7491 2927 7497
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3513 7531 3571 7537
rect 3513 7528 3525 7531
rect 3292 7500 3525 7528
rect 3292 7488 3298 7500
rect 3513 7497 3525 7500
rect 3559 7497 3571 7531
rect 3513 7491 3571 7497
rect 3878 7460 3884 7472
rect 2056 7432 2728 7460
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2700 7401 2728 7432
rect 3068 7432 3884 7460
rect 3068 7401 3096 7432
rect 3878 7420 3884 7432
rect 3936 7420 3942 7472
rect 4522 7420 4528 7472
rect 4580 7460 4586 7472
rect 4580 7432 6408 7460
rect 4580 7420 4586 7432
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 1912 7364 2145 7392
rect 1912 7352 1918 7364
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7361 3111 7395
rect 3053 7355 3111 7361
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 1302 7284 1308 7336
rect 1360 7324 1366 7336
rect 2608 7324 2636 7355
rect 3344 7324 3372 7355
rect 3786 7352 3792 7404
rect 3844 7352 3850 7404
rect 5810 7352 5816 7404
rect 5868 7352 5874 7404
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6380 7401 6408 7432
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 1360 7296 2636 7324
rect 2746 7296 3372 7324
rect 1360 7284 1366 7296
rect 1394 7216 1400 7268
rect 1452 7256 1458 7268
rect 1854 7256 1860 7268
rect 1452 7228 1860 7256
rect 1452 7216 1458 7228
rect 1854 7216 1860 7228
rect 1912 7216 1918 7268
rect 1946 7216 1952 7268
rect 2004 7256 2010 7268
rect 2409 7259 2467 7265
rect 2409 7256 2421 7259
rect 2004 7228 2421 7256
rect 2004 7216 2010 7228
rect 2409 7225 2421 7228
rect 2455 7225 2467 7259
rect 2409 7219 2467 7225
rect 1578 7148 1584 7200
rect 1636 7148 1642 7200
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2746 7188 2774 7296
rect 3237 7259 3295 7265
rect 3237 7225 3249 7259
rect 3283 7256 3295 7259
rect 4798 7256 4804 7268
rect 3283 7228 4804 7256
rect 3283 7225 3295 7228
rect 3237 7219 3295 7225
rect 4798 7216 4804 7228
rect 4856 7216 4862 7268
rect 4982 7216 4988 7268
rect 5040 7256 5046 7268
rect 5350 7256 5356 7268
rect 5040 7228 5356 7256
rect 5040 7216 5046 7228
rect 5350 7216 5356 7228
rect 5408 7256 5414 7268
rect 6549 7259 6607 7265
rect 6549 7256 6561 7259
rect 5408 7228 6561 7256
rect 5408 7216 5414 7228
rect 6549 7225 6561 7228
rect 6595 7225 6607 7259
rect 6549 7219 6607 7225
rect 2363 7160 2774 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 4672 7160 5089 7188
rect 4672 7148 4678 7160
rect 5077 7157 5089 7160
rect 5123 7157 5135 7191
rect 5077 7151 5135 7157
rect 5626 7148 5632 7200
rect 5684 7148 5690 7200
rect 6086 7148 6092 7200
rect 6144 7148 6150 7200
rect 1104 7098 6900 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 6900 7098
rect 1104 7024 6900 7046
rect 1854 6944 1860 6996
rect 1912 6944 1918 6996
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 3200 6956 4568 6984
rect 3200 6944 3206 6956
rect 1578 6876 1584 6928
rect 1636 6916 1642 6928
rect 3970 6916 3976 6928
rect 1636 6888 3976 6916
rect 1636 6876 1642 6888
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 4540 6925 4568 6956
rect 4525 6919 4583 6925
rect 4525 6885 4537 6919
rect 4571 6916 4583 6919
rect 5353 6919 5411 6925
rect 5353 6916 5365 6919
rect 4571 6888 5365 6916
rect 4571 6885 4583 6888
rect 4525 6879 4583 6885
rect 5353 6885 5365 6888
rect 5399 6885 5411 6919
rect 5353 6879 5411 6885
rect 1486 6808 1492 6860
rect 1544 6848 1550 6860
rect 1765 6851 1823 6857
rect 1765 6848 1777 6851
rect 1544 6820 1777 6848
rect 1544 6808 1550 6820
rect 1765 6817 1777 6820
rect 1811 6817 1823 6851
rect 4893 6851 4951 6857
rect 4893 6848 4905 6851
rect 1765 6811 1823 6817
rect 2148 6820 3740 6848
rect 1670 6740 1676 6792
rect 1728 6740 1734 6792
rect 1946 6740 1952 6792
rect 2004 6740 2010 6792
rect 2148 6712 2176 6820
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2498 6780 2504 6792
rect 2271 6752 2504 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 2590 6740 2596 6792
rect 2648 6740 2654 6792
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 1504 6684 2176 6712
rect 1504 6656 1532 6684
rect 2314 6672 2320 6724
rect 2372 6672 2378 6724
rect 2406 6672 2412 6724
rect 2464 6672 2470 6724
rect 2884 6712 2912 6743
rect 2958 6740 2964 6792
rect 3016 6740 3022 6792
rect 3142 6740 3148 6792
rect 3200 6740 3206 6792
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3418 6780 3424 6792
rect 3283 6752 3424 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 3602 6740 3608 6792
rect 3660 6740 3666 6792
rect 3712 6780 3740 6820
rect 3988 6820 4905 6848
rect 3988 6780 4016 6820
rect 4893 6817 4905 6820
rect 4939 6817 4951 6851
rect 4893 6811 4951 6817
rect 3712 6752 4016 6780
rect 4338 6740 4344 6792
rect 4396 6740 4402 6792
rect 4430 6740 4436 6792
rect 4488 6780 4494 6792
rect 4709 6783 4767 6789
rect 4709 6780 4721 6783
rect 4488 6752 4721 6780
rect 4488 6740 4494 6752
rect 4709 6749 4721 6752
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 2884 6684 3801 6712
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 4816 6712 4844 6743
rect 4982 6740 4988 6792
rect 5040 6740 5046 6792
rect 5258 6740 5264 6792
rect 5316 6740 5322 6792
rect 5442 6740 5448 6792
rect 5500 6780 5506 6792
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5500 6752 5917 6780
rect 5500 6740 5506 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 4028 6684 4844 6712
rect 5169 6715 5227 6721
rect 4028 6672 4034 6684
rect 5169 6681 5181 6715
rect 5215 6681 5227 6715
rect 5169 6675 5227 6681
rect 5629 6715 5687 6721
rect 5629 6681 5641 6715
rect 5675 6712 5687 6715
rect 5810 6712 5816 6724
rect 5675 6684 5816 6712
rect 5675 6681 5687 6684
rect 5629 6675 5687 6681
rect 1486 6604 1492 6656
rect 1544 6604 1550 6656
rect 2038 6604 2044 6656
rect 2096 6604 2102 6656
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 2685 6647 2743 6653
rect 2685 6644 2697 6647
rect 2188 6616 2697 6644
rect 2188 6604 2194 6616
rect 2685 6613 2697 6616
rect 2731 6613 2743 6647
rect 2685 6607 2743 6613
rect 3421 6647 3479 6653
rect 3421 6613 3433 6647
rect 3467 6644 3479 6647
rect 3878 6644 3884 6656
rect 3467 6616 3884 6644
rect 3467 6613 3479 6616
rect 3421 6607 3479 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5184 6644 5212 6675
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 4764 6616 5212 6644
rect 5537 6647 5595 6653
rect 4764 6604 4770 6616
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 6454 6644 6460 6656
rect 5583 6616 6460 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 6595 6616 6960 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 1104 6554 6900 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 6900 6554
rect 1104 6480 6900 6502
rect 1489 6443 1547 6449
rect 1489 6409 1501 6443
rect 1535 6440 1547 6443
rect 2406 6440 2412 6452
rect 1535 6412 2412 6440
rect 1535 6409 1547 6412
rect 1489 6403 1547 6409
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 3697 6443 3755 6449
rect 3697 6440 3709 6443
rect 2556 6412 3709 6440
rect 2556 6400 2562 6412
rect 3697 6409 3709 6412
rect 3743 6409 3755 6443
rect 3697 6403 3755 6409
rect 3878 6400 3884 6452
rect 3936 6440 3942 6452
rect 5534 6440 5540 6452
rect 3936 6412 5540 6440
rect 3936 6400 3942 6412
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 6454 6400 6460 6452
rect 6512 6400 6518 6452
rect 2130 6332 2136 6384
rect 2188 6332 2194 6384
rect 2774 6332 2780 6384
rect 2832 6332 2838 6384
rect 3602 6332 3608 6384
rect 3660 6332 3666 6384
rect 4614 6372 4620 6384
rect 4448 6344 4620 6372
rect 1486 6264 1492 6316
rect 1544 6264 1550 6316
rect 1578 6264 1584 6316
rect 1636 6264 1642 6316
rect 3620 6304 3648 6332
rect 4448 6313 4476 6344
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 4706 6332 4712 6384
rect 4764 6332 4770 6384
rect 4433 6307 4491 6313
rect 3620 6276 4384 6304
rect 1765 6239 1823 6245
rect 1765 6205 1777 6239
rect 1811 6205 1823 6239
rect 1765 6199 1823 6205
rect 1780 6168 1808 6199
rect 1854 6196 1860 6248
rect 1912 6196 1918 6248
rect 2498 6236 2504 6248
rect 1964 6208 2504 6236
rect 1964 6168 1992 6208
rect 2498 6196 2504 6208
rect 2556 6236 2562 6248
rect 2556 6208 3556 6236
rect 2556 6196 2562 6208
rect 1780 6140 1992 6168
rect 3528 6168 3556 6208
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 3660 6208 4261 6236
rect 3660 6196 3666 6208
rect 4249 6205 4261 6208
rect 4295 6205 4307 6239
rect 4356 6236 4384 6276
rect 4433 6273 4445 6307
rect 4479 6273 4491 6307
rect 6454 6304 6460 6316
rect 5842 6276 6460 6304
rect 4433 6267 4491 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 6932 6304 6960 6616
rect 6595 6276 6960 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 5442 6236 5448 6248
rect 4356 6208 5448 6236
rect 4249 6199 4307 6205
rect 5442 6196 5448 6208
rect 5500 6236 5506 6248
rect 6181 6239 6239 6245
rect 6181 6236 6193 6239
rect 5500 6208 6193 6236
rect 5500 6196 5506 6208
rect 6181 6205 6193 6208
rect 6227 6205 6239 6239
rect 6181 6199 6239 6205
rect 4430 6168 4436 6180
rect 3528 6140 4436 6168
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 1452 6072 3617 6100
rect 1452 6060 1458 6072
rect 3605 6069 3617 6072
rect 3651 6100 3663 6103
rect 4338 6100 4344 6112
rect 3651 6072 4344 6100
rect 3651 6069 3663 6072
rect 3605 6063 3663 6069
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 1104 6010 6900 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 6900 6010
rect 1104 5936 6900 5958
rect 1210 5856 1216 5908
rect 1268 5896 1274 5908
rect 1489 5899 1547 5905
rect 1489 5896 1501 5899
rect 1268 5868 1501 5896
rect 1268 5856 1274 5868
rect 1489 5865 1501 5868
rect 1535 5865 1547 5899
rect 1489 5859 1547 5865
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 2648 5868 3801 5896
rect 2648 5856 2654 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 3602 5788 3608 5840
rect 3660 5788 3666 5840
rect 4264 5800 4660 5828
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 4264 5760 4292 5800
rect 4632 5772 4660 5800
rect 1912 5732 4292 5760
rect 4433 5763 4491 5769
rect 1912 5720 1918 5732
rect 4433 5729 4445 5763
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 1673 5695 1731 5701
rect 1673 5692 1685 5695
rect 1452 5664 1685 5692
rect 1452 5652 1458 5664
rect 1673 5661 1685 5664
rect 1719 5661 1731 5695
rect 4448 5692 4476 5723
rect 4614 5720 4620 5772
rect 4672 5760 4678 5772
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 4672 5732 4813 5760
rect 4672 5720 4678 5732
rect 4801 5729 4813 5732
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 4706 5692 4712 5704
rect 4448 5664 4712 5692
rect 1673 5655 1731 5661
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 2038 5584 2044 5636
rect 2096 5624 2102 5636
rect 2133 5627 2191 5633
rect 2133 5624 2145 5627
rect 2096 5596 2145 5624
rect 2096 5584 2102 5596
rect 2133 5593 2145 5596
rect 2179 5593 2191 5627
rect 2133 5587 2191 5593
rect 3142 5584 3148 5636
rect 3200 5584 3206 5636
rect 4157 5627 4215 5633
rect 4157 5593 4169 5627
rect 4203 5624 4215 5627
rect 4614 5624 4620 5636
rect 4203 5596 4620 5624
rect 4203 5593 4215 5596
rect 4157 5587 4215 5593
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 5077 5627 5135 5633
rect 5077 5593 5089 5627
rect 5123 5624 5135 5627
rect 5350 5624 5356 5636
rect 5123 5596 5356 5624
rect 5123 5593 5135 5596
rect 5077 5587 5135 5593
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 6638 5624 6644 5636
rect 6302 5596 6644 5624
rect 6638 5584 6644 5596
rect 6696 5584 6702 5636
rect 3418 5516 3424 5568
rect 3476 5556 3482 5568
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 3476 5528 4261 5556
rect 3476 5516 3482 5528
rect 4249 5525 4261 5528
rect 4295 5556 4307 5559
rect 4706 5556 4712 5568
rect 4295 5528 4712 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4706 5516 4712 5528
rect 4764 5556 4770 5568
rect 5258 5556 5264 5568
rect 4764 5528 5264 5556
rect 4764 5516 4770 5528
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 6546 5516 6552 5568
rect 6604 5516 6610 5568
rect 1104 5466 6900 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 6900 5466
rect 1104 5392 6900 5414
rect 1302 5312 1308 5364
rect 1360 5352 1366 5364
rect 1489 5355 1547 5361
rect 1489 5352 1501 5355
rect 1360 5324 1501 5352
rect 1360 5312 1366 5324
rect 1489 5321 1501 5324
rect 1535 5321 1547 5355
rect 1489 5315 1547 5321
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 1765 5355 1823 5361
rect 1765 5352 1777 5355
rect 1728 5324 1777 5352
rect 1728 5312 1734 5324
rect 1765 5321 1777 5324
rect 1811 5321 1823 5355
rect 1765 5315 1823 5321
rect 1946 5312 1952 5364
rect 2004 5352 2010 5364
rect 2041 5355 2099 5361
rect 2041 5352 2053 5355
rect 2004 5324 2053 5352
rect 2004 5312 2010 5324
rect 2041 5321 2053 5324
rect 2087 5321 2099 5355
rect 2041 5315 2099 5321
rect 2498 5312 2504 5364
rect 2556 5312 2562 5364
rect 2774 5312 2780 5364
rect 2832 5312 2838 5364
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3142 5352 3148 5364
rect 3099 5324 3148 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3142 5312 3148 5324
rect 3200 5312 3206 5364
rect 5445 5355 5503 5361
rect 5445 5321 5457 5355
rect 5491 5352 5503 5355
rect 5902 5352 5908 5364
rect 5491 5324 5908 5352
rect 5491 5321 5503 5324
rect 5445 5315 5503 5321
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 3602 5284 3608 5296
rect 1688 5256 3608 5284
rect 1688 5225 1716 5256
rect 3602 5244 3608 5256
rect 3660 5244 3666 5296
rect 4798 5244 4804 5296
rect 4856 5284 4862 5296
rect 5350 5284 5356 5296
rect 4856 5256 5356 5284
rect 4856 5244 4862 5256
rect 5350 5244 5356 5256
rect 5408 5284 5414 5296
rect 5408 5256 6592 5284
rect 5408 5244 5414 5256
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 1762 5176 1768 5228
rect 1820 5216 1826 5228
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1820 5188 1961 5216
rect 1820 5176 1826 5188
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2222 5176 2228 5228
rect 2280 5176 2286 5228
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 3145 5219 3203 5225
rect 3145 5216 3157 5219
rect 2915 5188 3157 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 3145 5185 3157 5188
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 1210 5108 1216 5160
rect 1268 5148 1274 5160
rect 2332 5148 2360 5179
rect 1268 5120 2360 5148
rect 3160 5148 3188 5179
rect 3234 5176 3240 5228
rect 3292 5176 3298 5228
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5442 5216 5448 5228
rect 5307 5188 5448 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 6564 5225 6592 5256
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 3602 5148 3608 5160
rect 3160 5120 3608 5148
rect 1268 5108 1274 5120
rect 3602 5108 3608 5120
rect 3660 5148 3666 5160
rect 5626 5148 5632 5160
rect 3660 5120 5632 5148
rect 3660 5108 3666 5120
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 6178 5108 6184 5160
rect 6236 5108 6242 5160
rect 3786 4972 3792 5024
rect 3844 5012 3850 5024
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 3844 4984 4537 5012
rect 3844 4972 3850 4984
rect 4525 4981 4537 4984
rect 4571 4981 4583 5015
rect 4525 4975 4583 4981
rect 5534 4972 5540 5024
rect 5592 4972 5598 5024
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 5868 4984 6469 5012
rect 5868 4972 5874 4984
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6457 4975 6515 4981
rect 1104 4922 6900 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 6900 4922
rect 1104 4848 6900 4870
rect 4246 4808 4252 4820
rect 3160 4780 4252 4808
rect 3160 4613 3188 4780
rect 4246 4768 4252 4780
rect 4304 4808 4310 4820
rect 4614 4808 4620 4820
rect 4304 4780 4620 4808
rect 4304 4768 4310 4780
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 4154 4700 4160 4752
rect 4212 4700 4218 4752
rect 4341 4743 4399 4749
rect 4341 4709 4353 4743
rect 4387 4740 4399 4743
rect 4706 4740 4712 4752
rect 4387 4712 4712 4740
rect 4387 4709 4399 4712
rect 4341 4703 4399 4709
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 5626 4700 5632 4752
rect 5684 4700 5690 4752
rect 5905 4675 5963 4681
rect 5905 4672 5917 4675
rect 3620 4644 5917 4672
rect 3620 4613 3648 4644
rect 5905 4641 5917 4644
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4573 3663 4607
rect 3605 4567 3663 4573
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 3752 4576 3801 4604
rect 3752 4564 3758 4576
rect 3789 4573 3801 4576
rect 3835 4604 3847 4607
rect 4525 4607 4583 4613
rect 4525 4604 4537 4607
rect 3835 4576 4537 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 4525 4573 4537 4576
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 4798 4604 4804 4616
rect 4755 4576 4804 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 3326 4496 3332 4548
rect 3384 4496 3390 4548
rect 4154 4496 4160 4548
rect 4212 4536 4218 4548
rect 4724 4536 4752 4567
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4573 5043 4607
rect 4985 4567 5043 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4604 5503 4607
rect 5534 4604 5540 4616
rect 5491 4576 5540 4604
rect 5491 4573 5503 4576
rect 5445 4567 5503 4573
rect 4212 4508 4752 4536
rect 5000 4536 5028 4567
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6236 4576 6469 4604
rect 6236 4564 6242 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 6196 4536 6224 4564
rect 5000 4508 6224 4536
rect 4212 4496 4218 4508
rect 2958 4428 2964 4480
rect 3016 4428 3022 4480
rect 3513 4471 3571 4477
rect 3513 4437 3525 4471
rect 3559 4468 3571 4471
rect 3878 4468 3884 4480
rect 3559 4440 3884 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 5169 4471 5227 4477
rect 5169 4437 5181 4471
rect 5215 4468 5227 4471
rect 5258 4468 5264 4480
rect 5215 4440 5264 4468
rect 5215 4437 5227 4440
rect 5169 4431 5227 4437
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 1104 4378 6900 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 6900 4378
rect 1104 4304 6900 4326
rect 3326 4224 3332 4276
rect 3384 4264 3390 4276
rect 3421 4267 3479 4273
rect 3421 4264 3433 4267
rect 3384 4236 3433 4264
rect 3384 4224 3390 4236
rect 3421 4233 3433 4236
rect 3467 4233 3479 4267
rect 4246 4264 4252 4276
rect 3421 4227 3479 4233
rect 3528 4236 4252 4264
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2731 4100 2973 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2961 4097 2973 4100
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 3053 4131 3111 4137
rect 3053 4097 3065 4131
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 1670 4020 1676 4072
rect 1728 4060 1734 4072
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 1728 4032 2053 4060
rect 1728 4020 1734 4032
rect 2041 4029 2053 4032
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 3068 4060 3096 4091
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 3200 4100 3249 4128
rect 3200 4088 3206 4100
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 3528 4128 3556 4236
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 5626 4224 5632 4276
rect 5684 4264 5690 4276
rect 5684 4236 6408 4264
rect 5684 4224 5690 4236
rect 3878 4156 3884 4208
rect 3936 4156 3942 4208
rect 6270 4196 6276 4208
rect 5934 4168 6276 4196
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 3375 4100 3556 4128
rect 3605 4131 3663 4137
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 3605 4097 3617 4131
rect 3651 4128 3663 4131
rect 3694 4128 3700 4140
rect 3651 4100 3700 4128
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 3970 4128 3976 4140
rect 3804 4100 3976 4128
rect 3804 4069 3832 4100
rect 3970 4088 3976 4100
rect 4028 4128 4034 4140
rect 4065 4131 4123 4137
rect 4065 4128 4077 4131
rect 4028 4100 4077 4128
rect 4028 4088 4034 4100
rect 4065 4097 4077 4100
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 6380 4137 6408 4236
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 3789 4063 3847 4069
rect 3789 4060 3801 4063
rect 2924 4032 3801 4060
rect 2924 4020 2930 4032
rect 3789 4029 3801 4032
rect 3835 4029 3847 4063
rect 3789 4023 3847 4029
rect 4430 4020 4436 4072
rect 4488 4020 4494 4072
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 4540 4032 4721 4060
rect 3142 3952 3148 4004
rect 3200 3992 3206 4004
rect 4157 3995 4215 4001
rect 4157 3992 4169 3995
rect 3200 3964 4169 3992
rect 3200 3952 3206 3964
rect 4157 3961 4169 3964
rect 4203 3961 4215 3995
rect 4157 3955 4215 3961
rect 4341 3995 4399 4001
rect 4341 3961 4353 3995
rect 4387 3992 4399 3995
rect 4540 3992 4568 4032
rect 4709 4029 4721 4032
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 4387 3964 4568 3992
rect 6380 3992 6408 4091
rect 6454 4088 6460 4140
rect 6512 4088 6518 4140
rect 6454 3992 6460 4004
rect 6380 3964 6460 3992
rect 4387 3961 4399 3964
rect 4341 3955 4399 3961
rect 2777 3927 2835 3933
rect 2777 3893 2789 3927
rect 2823 3924 2835 3927
rect 3050 3924 3056 3936
rect 2823 3896 3056 3924
rect 2823 3893 2835 3896
rect 2777 3887 2835 3893
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 4172 3924 4200 3955
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 4706 3924 4712 3936
rect 4172 3896 4712 3924
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 6178 3924 6184 3936
rect 5776 3896 6184 3924
rect 5776 3884 5782 3896
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 1104 3834 6900 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 6900 3834
rect 1104 3760 6900 3782
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 3694 3720 3700 3732
rect 3651 3692 3700 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 3694 3680 3700 3692
rect 3752 3720 3758 3732
rect 4062 3720 4068 3732
rect 3752 3692 4068 3720
rect 3752 3680 3758 3692
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4430 3680 4436 3732
rect 4488 3720 4494 3732
rect 4706 3720 4712 3732
rect 4488 3692 4712 3720
rect 4488 3680 4494 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 6362 3680 6368 3732
rect 6420 3680 6426 3732
rect 842 3612 848 3664
rect 900 3652 906 3664
rect 1489 3655 1547 3661
rect 1489 3652 1501 3655
rect 900 3624 1501 3652
rect 900 3612 906 3624
rect 1489 3621 1501 3624
rect 1535 3621 1547 3655
rect 1489 3615 1547 3621
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3584 1915 3587
rect 4341 3587 4399 3593
rect 4341 3584 4353 3587
rect 1903 3556 4353 3584
rect 1903 3553 1915 3556
rect 1857 3547 1915 3553
rect 4341 3553 4353 3556
rect 4387 3584 4399 3587
rect 4614 3584 4620 3596
rect 4387 3556 4620 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 1670 3476 1676 3528
rect 1728 3476 1734 3528
rect 3694 3476 3700 3528
rect 3752 3516 3758 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3752 3488 3801 3516
rect 3752 3476 3758 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 3970 3476 3976 3528
rect 4028 3476 4034 3528
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 2133 3451 2191 3457
rect 2133 3417 2145 3451
rect 2179 3417 2191 3451
rect 3510 3448 3516 3460
rect 3358 3420 3516 3448
rect 2133 3411 2191 3417
rect 2148 3380 2176 3411
rect 3510 3408 3516 3420
rect 3568 3408 3574 3460
rect 3602 3408 3608 3460
rect 3660 3448 3666 3460
rect 4080 3448 4108 3479
rect 6546 3476 6552 3528
rect 6604 3476 6610 3528
rect 3660 3420 4108 3448
rect 3660 3408 3666 3420
rect 4522 3408 4528 3460
rect 4580 3448 4586 3460
rect 4617 3451 4675 3457
rect 4617 3448 4629 3451
rect 4580 3420 4629 3448
rect 4580 3408 4586 3420
rect 4617 3417 4629 3420
rect 4663 3417 4675 3451
rect 4617 3411 4675 3417
rect 4724 3420 5106 3448
rect 2958 3380 2964 3392
rect 2148 3352 2964 3380
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 3878 3340 3884 3392
rect 3936 3340 3942 3392
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4724 3380 4752 3420
rect 4203 3352 4752 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 6086 3340 6092 3392
rect 6144 3340 6150 3392
rect 1104 3290 6900 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 6900 3290
rect 1104 3216 6900 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 1670 3176 1676 3188
rect 1627 3148 1676 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 3510 3136 3516 3188
rect 3568 3136 3574 3188
rect 3970 3136 3976 3188
rect 4028 3176 4034 3188
rect 4028 3148 4476 3176
rect 4028 3136 4034 3148
rect 2958 3108 2964 3120
rect 2622 3080 2964 3108
rect 2958 3068 2964 3080
rect 3016 3068 3022 3120
rect 3050 3068 3056 3120
rect 3108 3068 3114 3120
rect 3878 3068 3884 3120
rect 3936 3108 3942 3120
rect 4448 3108 4476 3148
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 4580 3148 4905 3176
rect 4580 3136 4586 3148
rect 4893 3145 4905 3148
rect 4939 3145 4951 3179
rect 4893 3139 4951 3145
rect 6457 3179 6515 3185
rect 6457 3145 6469 3179
rect 6503 3176 6515 3179
rect 6638 3176 6644 3188
rect 6503 3148 6644 3176
rect 6503 3145 6515 3148
rect 6457 3139 6515 3145
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 5810 3108 5816 3120
rect 3936 3080 4384 3108
rect 4448 3080 5816 3108
rect 3936 3068 3942 3080
rect 3602 3000 3608 3052
rect 3660 3000 3666 3052
rect 4062 3000 4068 3052
rect 4120 3000 4126 3052
rect 4356 3049 4384 3080
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 4430 3000 4436 3052
rect 4488 3000 4494 3052
rect 4632 3049 4660 3080
rect 5810 3068 5816 3080
rect 5868 3068 5874 3120
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 6086 3040 6092 3052
rect 5399 3012 6092 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 3344 2836 3372 2935
rect 3694 2932 3700 2984
rect 3752 2932 3758 2984
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2972 4031 2975
rect 4724 2972 4752 3003
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 6454 3040 6460 3052
rect 6411 3012 6460 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 5445 2975 5503 2981
rect 5445 2972 5457 2975
rect 4019 2944 4660 2972
rect 4724 2944 5457 2972
rect 4019 2941 4031 2944
rect 3973 2935 4031 2941
rect 4632 2904 4660 2944
rect 5445 2941 5457 2944
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 5626 2904 5632 2916
rect 4632 2876 5632 2904
rect 5626 2864 5632 2876
rect 5684 2864 5690 2916
rect 4614 2836 4620 2848
rect 3344 2808 4620 2836
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 5166 2796 5172 2848
rect 5224 2796 5230 2848
rect 1104 2746 6900 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 6900 2746
rect 1104 2672 6900 2694
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3237 2635 3295 2641
rect 3237 2632 3249 2635
rect 3016 2604 3249 2632
rect 3016 2592 3022 2604
rect 3237 2601 3249 2604
rect 3283 2601 3295 2635
rect 3237 2595 3295 2601
rect 4614 2592 4620 2644
rect 4672 2632 4678 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 4672 2604 5089 2632
rect 4672 2592 4678 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 5626 2592 5632 2644
rect 5684 2592 5690 2644
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 6178 2632 6184 2644
rect 6135 2604 6184 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 6270 2592 6276 2644
rect 6328 2632 6334 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 6328 2604 6469 2632
rect 6328 2592 6334 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 3605 2567 3663 2573
rect 3605 2533 3617 2567
rect 3651 2533 3663 2567
rect 3605 2527 3663 2533
rect 3510 2496 3516 2508
rect 3344 2468 3516 2496
rect 3344 2437 3372 2468
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 3620 2496 3648 2527
rect 3620 2468 5948 2496
rect 3329 2431 3387 2437
rect 3329 2397 3341 2431
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 3436 2360 3464 2391
rect 3786 2388 3792 2440
rect 3844 2388 3850 2440
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 5920 2437 5948 2468
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 4580 2400 5825 2428
rect 4580 2388 4586 2400
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 6454 2428 6460 2440
rect 6411 2400 6460 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 5718 2360 5724 2372
rect 3436 2332 5724 2360
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 1104 2202 6900 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 6900 2202
rect 1104 2128 6900 2150
<< via1 >>
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1952 7420 2004 7472
rect 2596 7488 2648 7540
rect 3240 7488 3292 7540
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 3884 7420 3936 7472
rect 4528 7420 4580 7472
rect 1860 7352 1912 7361
rect 1308 7284 1360 7336
rect 3792 7395 3844 7404
rect 3792 7361 3801 7395
rect 3801 7361 3835 7395
rect 3835 7361 3844 7395
rect 3792 7352 3844 7361
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 1400 7216 1452 7268
rect 1860 7216 1912 7268
rect 1952 7216 2004 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 4804 7216 4856 7268
rect 4988 7216 5040 7268
rect 5356 7216 5408 7268
rect 4620 7148 4672 7200
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 6092 7191 6144 7200
rect 6092 7157 6101 7191
rect 6101 7157 6135 7191
rect 6135 7157 6144 7191
rect 6092 7148 6144 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1860 6987 1912 6996
rect 1860 6953 1869 6987
rect 1869 6953 1903 6987
rect 1903 6953 1912 6987
rect 1860 6944 1912 6953
rect 3148 6944 3200 6996
rect 1584 6876 1636 6928
rect 3976 6876 4028 6928
rect 1492 6808 1544 6860
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 2504 6740 2556 6792
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 2320 6715 2372 6724
rect 2320 6681 2329 6715
rect 2329 6681 2363 6715
rect 2363 6681 2372 6715
rect 2320 6672 2372 6681
rect 2412 6715 2464 6724
rect 2412 6681 2421 6715
rect 2421 6681 2455 6715
rect 2455 6681 2464 6715
rect 2412 6672 2464 6681
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 3424 6740 3476 6792
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 4436 6740 4488 6792
rect 3976 6672 4028 6724
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 5448 6740 5500 6792
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 2136 6604 2188 6656
rect 3884 6604 3936 6656
rect 4712 6604 4764 6656
rect 5816 6672 5868 6724
rect 6460 6604 6512 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2412 6400 2464 6452
rect 2504 6400 2556 6452
rect 3884 6400 3936 6452
rect 5540 6400 5592 6452
rect 6460 6443 6512 6452
rect 6460 6409 6469 6443
rect 6469 6409 6503 6443
rect 6503 6409 6512 6443
rect 6460 6400 6512 6409
rect 2136 6375 2188 6384
rect 2136 6341 2145 6375
rect 2145 6341 2179 6375
rect 2179 6341 2188 6375
rect 2136 6332 2188 6341
rect 2780 6332 2832 6384
rect 3608 6332 3660 6384
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 1492 6264 1544 6273
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 4620 6332 4672 6384
rect 4712 6375 4764 6384
rect 4712 6341 4721 6375
rect 4721 6341 4755 6375
rect 4755 6341 4764 6375
rect 4712 6332 4764 6341
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 2504 6196 2556 6248
rect 3608 6196 3660 6248
rect 6460 6264 6512 6316
rect 5448 6196 5500 6248
rect 4436 6128 4488 6180
rect 1400 6060 1452 6112
rect 4344 6060 4396 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 1216 5856 1268 5908
rect 2596 5856 2648 5908
rect 3608 5831 3660 5840
rect 3608 5797 3617 5831
rect 3617 5797 3651 5831
rect 3651 5797 3660 5831
rect 3608 5788 3660 5797
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 1400 5652 1452 5704
rect 4620 5720 4672 5772
rect 4712 5652 4764 5704
rect 2044 5584 2096 5636
rect 3148 5584 3200 5636
rect 4620 5584 4672 5636
rect 5356 5584 5408 5636
rect 6644 5584 6696 5636
rect 3424 5516 3476 5568
rect 4712 5516 4764 5568
rect 5264 5516 5316 5568
rect 6552 5559 6604 5568
rect 6552 5525 6561 5559
rect 6561 5525 6595 5559
rect 6595 5525 6604 5559
rect 6552 5516 6604 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 1308 5312 1360 5364
rect 1676 5312 1728 5364
rect 1952 5312 2004 5364
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 3148 5312 3200 5364
rect 5908 5312 5960 5364
rect 3608 5244 3660 5296
rect 4804 5244 4856 5296
rect 5356 5244 5408 5296
rect 1768 5176 1820 5228
rect 2228 5219 2280 5228
rect 2228 5185 2237 5219
rect 2237 5185 2271 5219
rect 2271 5185 2280 5219
rect 2228 5176 2280 5185
rect 1216 5108 1268 5160
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 5448 5176 5500 5228
rect 3608 5108 3660 5160
rect 5632 5108 5684 5160
rect 6184 5151 6236 5160
rect 6184 5117 6193 5151
rect 6193 5117 6227 5151
rect 6227 5117 6236 5151
rect 6184 5108 6236 5117
rect 3792 4972 3844 5024
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 5816 4972 5868 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 4252 4811 4304 4820
rect 4252 4777 4261 4811
rect 4261 4777 4295 4811
rect 4295 4777 4304 4811
rect 4252 4768 4304 4777
rect 4620 4768 4672 4820
rect 4160 4743 4212 4752
rect 4160 4709 4169 4743
rect 4169 4709 4203 4743
rect 4203 4709 4212 4743
rect 4160 4700 4212 4709
rect 4712 4700 4764 4752
rect 5632 4743 5684 4752
rect 5632 4709 5641 4743
rect 5641 4709 5675 4743
rect 5675 4709 5684 4743
rect 5632 4700 5684 4709
rect 3700 4564 3752 4616
rect 3332 4539 3384 4548
rect 3332 4505 3341 4539
rect 3341 4505 3375 4539
rect 3375 4505 3384 4539
rect 3332 4496 3384 4505
rect 4160 4496 4212 4548
rect 4804 4564 4856 4616
rect 5540 4564 5592 4616
rect 6184 4564 6236 4616
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 3884 4428 3936 4480
rect 5264 4428 5316 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 3332 4224 3384 4276
rect 1676 4020 1728 4072
rect 2872 4020 2924 4072
rect 3148 4088 3200 4140
rect 4252 4224 4304 4276
rect 5632 4224 5684 4276
rect 3884 4199 3936 4208
rect 3884 4165 3893 4199
rect 3893 4165 3927 4199
rect 3927 4165 3936 4199
rect 3884 4156 3936 4165
rect 6276 4156 6328 4208
rect 3700 4088 3752 4140
rect 3976 4088 4028 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 4436 4063 4488 4072
rect 4436 4029 4445 4063
rect 4445 4029 4479 4063
rect 4479 4029 4488 4063
rect 4436 4020 4488 4029
rect 3148 3952 3200 4004
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 3056 3884 3108 3936
rect 6460 3952 6512 4004
rect 4712 3884 4764 3936
rect 5724 3884 5776 3936
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 3700 3680 3752 3732
rect 4068 3680 4120 3732
rect 4436 3680 4488 3732
rect 4712 3680 4764 3732
rect 6368 3723 6420 3732
rect 6368 3689 6377 3723
rect 6377 3689 6411 3723
rect 6411 3689 6420 3723
rect 6368 3680 6420 3689
rect 848 3612 900 3664
rect 4620 3544 4672 3596
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 3700 3476 3752 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 3516 3408 3568 3460
rect 3608 3408 3660 3460
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 4528 3408 4580 3460
rect 2964 3340 3016 3392
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 6092 3383 6144 3392
rect 6092 3349 6101 3383
rect 6101 3349 6135 3383
rect 6135 3349 6144 3383
rect 6092 3340 6144 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1676 3136 1728 3188
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 3976 3136 4028 3188
rect 2964 3068 3016 3120
rect 3056 3111 3108 3120
rect 3056 3077 3065 3111
rect 3065 3077 3099 3111
rect 3099 3077 3108 3111
rect 3056 3068 3108 3077
rect 3884 3068 3936 3120
rect 4528 3136 4580 3188
rect 6644 3136 6696 3188
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 4068 3043 4120 3052
rect 4068 3009 4077 3043
rect 4077 3009 4111 3043
rect 4111 3009 4120 3043
rect 4068 3000 4120 3009
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 5816 3068 5868 3120
rect 6092 3043 6144 3052
rect 3700 2975 3752 2984
rect 3700 2941 3709 2975
rect 3709 2941 3743 2975
rect 3743 2941 3752 2975
rect 3700 2932 3752 2941
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 6460 3000 6512 3052
rect 5632 2864 5684 2916
rect 4620 2796 4672 2848
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 5172 2796 5224 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 2964 2592 3016 2644
rect 4620 2592 4672 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 6184 2592 6236 2644
rect 6276 2592 6328 2644
rect 3516 2456 3568 2508
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 4528 2388 4580 2440
rect 6460 2388 6512 2440
rect 5724 2320 5776 2372
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 1950 9411 2006 10211
rect 2594 9411 2650 10211
rect 3238 9411 3294 10211
rect 3882 9411 3938 10211
rect 4526 9411 4582 10211
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1320 7342 1348 8191
rect 1766 7576 1822 7585
rect 1766 7511 1822 7520
rect 1308 7336 1360 7342
rect 1308 7278 1360 7284
rect 1400 7268 1452 7274
rect 1400 7210 1452 7216
rect 1214 6216 1270 6225
rect 1214 6151 1270 6160
rect 1228 5914 1256 6151
rect 1412 6118 1440 7210
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6934 1624 7142
rect 1584 6928 1636 6934
rect 1584 6870 1636 6876
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1504 6769 1532 6802
rect 1490 6760 1546 6769
rect 1490 6695 1546 6704
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6322 1532 6598
rect 1596 6322 1624 6870
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1216 5908 1268 5914
rect 1216 5850 1268 5856
rect 1412 5710 1440 6054
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1306 5536 1362 5545
rect 1306 5471 1362 5480
rect 1320 5370 1348 5471
rect 1688 5370 1716 6734
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1780 5234 1808 7511
rect 1964 7478 1992 9411
rect 2226 8936 2282 8945
rect 2226 8871 2282 8880
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1872 7274 1900 7346
rect 1860 7268 1912 7274
rect 1860 7210 1912 7216
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1872 6338 1900 6938
rect 1964 6798 1992 7210
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1872 6310 1992 6338
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1872 5778 1900 6190
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1964 5370 1992 6310
rect 2056 5642 2084 6598
rect 2148 6390 2176 6598
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2044 5636 2096 5642
rect 2044 5578 2096 5584
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 2240 5234 2268 8871
rect 2608 7546 2636 9411
rect 3252 7546 3280 9411
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3896 7478 3924 9411
rect 4540 7478 4568 9411
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3160 6798 3188 6938
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2332 6633 2360 6666
rect 2318 6624 2374 6633
rect 2318 6559 2374 6568
rect 2424 6458 2452 6666
rect 2516 6458 2544 6734
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2516 5370 2544 6190
rect 2608 5914 2636 6734
rect 2976 6633 3004 6734
rect 2962 6624 3018 6633
rect 2884 6582 2962 6610
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2792 5370 2820 6326
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 1216 5160 1268 5166
rect 1216 5102 1268 5108
rect 1228 4865 1256 5102
rect 1214 4856 1270 4865
rect 1214 4791 1270 4800
rect 2884 4078 2912 6582
rect 2962 6559 3018 6568
rect 3160 5896 3188 6734
rect 3068 5868 3188 5896
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 848 3664 900 3670
rect 846 3632 848 3641
rect 900 3632 902 3641
rect 846 3567 902 3576
rect 1688 3534 1716 4014
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1688 3194 1716 3470
rect 2976 3398 3004 4422
rect 3068 4162 3096 5868
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3160 5370 3188 5578
rect 3436 5574 3464 6734
rect 3620 6390 3648 6734
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5846 3648 6190
rect 3608 5840 3660 5846
rect 3608 5782 3660 5788
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3620 5302 3648 5782
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3252 4185 3280 5170
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3332 4548 3384 4554
rect 3332 4490 3384 4496
rect 3344 4282 3372 4490
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3238 4176 3294 4185
rect 3068 4146 3188 4162
rect 3068 4140 3200 4146
rect 3068 4134 3148 4140
rect 3238 4111 3294 4120
rect 3148 4082 3200 4088
rect 3160 4010 3188 4082
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 3068 3126 3096 3878
rect 3620 3466 3648 5102
rect 3804 5030 3832 7346
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3988 6730 4016 6870
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6458 3924 6598
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 4356 6118 4384 6734
rect 4448 6186 4476 6734
rect 4632 6390 4660 7142
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4724 6390 4752 6598
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5778 4660 6326
rect 4816 5794 4844 7210
rect 5000 6798 5028 7210
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4724 5766 4844 5794
rect 4724 5710 4752 5766
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3712 4146 3740 4558
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3712 3738 3740 4082
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3516 3460 3568 3466
rect 3516 3402 3568 3408
rect 3608 3460 3660 3466
rect 3608 3402 3660 3408
rect 3528 3194 3556 3402
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 2976 2650 3004 3062
rect 3620 3058 3648 3402
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3620 2530 3648 2994
rect 3712 2990 3740 3470
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3528 2514 3648 2530
rect 3516 2508 3648 2514
rect 3568 2502 3648 2508
rect 3516 2450 3568 2456
rect 3804 2446 3832 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4826 4660 5578
rect 5276 5574 5304 6734
rect 5368 5642 5396 7210
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5448 6792 5500 6798
rect 5644 6769 5672 7142
rect 5828 6905 5856 7346
rect 5814 6896 5870 6905
rect 5814 6831 5870 6840
rect 5448 6734 5500 6740
rect 5630 6760 5686 6769
rect 5460 6254 5488 6734
rect 5630 6695 5686 6704
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 6248 5500 6254
rect 5552 6225 5580 6394
rect 5448 6190 5500 6196
rect 5538 6216 5594 6225
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 4172 4554 4200 4694
rect 4160 4548 4212 4554
rect 4160 4490 4212 4496
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3896 4214 3924 4422
rect 4264 4282 4292 4762
rect 4724 4758 4752 5510
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5368 5302 5396 5578
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4816 4622 4844 5238
rect 5460 5234 5488 6190
rect 5538 6151 5594 6160
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4622 5580 4966
rect 5644 4758 5672 5102
rect 5828 5030 5856 6666
rect 5920 5370 5948 7346
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 6905 6132 7142
rect 6090 6896 6146 6905
rect 6090 6831 6146 6840
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6472 6458 6500 6598
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6366 5536 6422 5545
rect 6366 5471 6422 5480
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 4264 4146 4292 4218
rect 5276 4185 5304 4422
rect 5644 4282 5672 4694
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5262 4176 5318 4185
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4252 4140 4304 4146
rect 5262 4111 5318 4120
rect 4252 4082 4304 4088
rect 3988 3534 4016 4082
rect 4436 4072 4488 4078
rect 4488 4020 4660 4026
rect 4436 4014 4660 4020
rect 4448 3998 4660 4014
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3126 3924 3334
rect 3988 3194 4016 3470
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 4080 3058 4108 3674
rect 4448 3058 4476 3674
rect 4632 3602 4660 3998
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 4724 3738 4752 3878
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 4540 3194 4568 3402
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4632 2854 4660 3538
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 4620 2848 4672 2854
rect 5172 2848 5224 2854
rect 4620 2790 4672 2796
rect 5170 2816 5172 2825
rect 5224 2816 5226 2825
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 2790
rect 5170 2751 5226 2760
rect 5644 2650 5672 2858
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4540 800 4568 2382
rect 5736 2378 5764 3878
rect 5828 3126 5856 4966
rect 6196 4865 6224 5102
rect 6182 4856 6238 4865
rect 6182 4791 6238 4800
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6196 3942 6224 4558
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6182 3496 6238 3505
rect 6182 3431 6238 3440
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 6104 3058 6132 3334
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6196 2650 6224 3431
rect 6288 2650 6316 4150
rect 6380 3738 6408 5471
rect 6472 4146 6500 6258
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6472 3058 6500 3946
rect 6564 3534 6592 5510
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6656 3194 6684 5578
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6472 2446 6500 2994
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 4526 0 4582 800
<< via2 >>
rect 1306 8200 1362 8256
rect 1766 7520 1822 7576
rect 1214 6160 1270 6216
rect 1490 6704 1546 6760
rect 1306 5480 1362 5536
rect 2226 8880 2282 8936
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 2318 6568 2374 6624
rect 1214 4800 1270 4856
rect 2962 6568 3018 6624
rect 846 3612 848 3632
rect 848 3612 900 3632
rect 900 3612 902 3632
rect 846 3576 902 3612
rect 3238 4120 3294 4176
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 5814 6840 5870 6896
rect 5630 6704 5686 6760
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 5538 6160 5594 6216
rect 6090 6840 6146 6896
rect 6366 5480 6422 5536
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 5262 4120 5318 4176
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 5170 2796 5172 2816
rect 5172 2796 5224 2816
rect 5224 2796 5226 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5170 2760 5226 2796
rect 6182 4800 6238 4856
rect 6182 3440 6238 3496
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 0 8938 800 8968
rect 2221 8938 2287 8941
rect 0 8936 2287 8938
rect 0 8880 2226 8936
rect 2282 8880 2287 8936
rect 0 8878 2287 8880
rect 0 8848 800 8878
rect 2221 8875 2287 8878
rect 0 8258 800 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 0 8168 800 8198
rect 1301 8195 1367 8198
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 1761 7578 1827 7581
rect 0 7576 1827 7578
rect 0 7520 1766 7576
rect 1822 7520 1827 7576
rect 0 7518 1827 7520
rect 0 7488 800 7518
rect 1761 7515 1827 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 5809 6898 5875 6901
rect 0 6896 5875 6898
rect 0 6840 5814 6896
rect 5870 6840 5875 6896
rect 0 6838 5875 6840
rect 0 6808 800 6838
rect 5809 6835 5875 6838
rect 6085 6898 6151 6901
rect 7267 6898 8067 6928
rect 6085 6896 8067 6898
rect 6085 6840 6090 6896
rect 6146 6840 8067 6896
rect 6085 6838 8067 6840
rect 6085 6835 6151 6838
rect 7267 6808 8067 6838
rect 1485 6762 1551 6765
rect 5625 6762 5691 6765
rect 1485 6760 5691 6762
rect 1485 6704 1490 6760
rect 1546 6704 5630 6760
rect 5686 6704 5691 6760
rect 1485 6702 5691 6704
rect 1485 6699 1551 6702
rect 5625 6699 5691 6702
rect 2313 6626 2379 6629
rect 2957 6626 3023 6629
rect 2313 6624 3023 6626
rect 2313 6568 2318 6624
rect 2374 6568 2962 6624
rect 3018 6568 3023 6624
rect 2313 6566 3023 6568
rect 2313 6563 2379 6566
rect 2957 6563 3023 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 0 6218 800 6248
rect 1209 6218 1275 6221
rect 0 6216 1275 6218
rect 0 6160 1214 6216
rect 1270 6160 1275 6216
rect 0 6158 1275 6160
rect 0 6128 800 6158
rect 1209 6155 1275 6158
rect 5533 6218 5599 6221
rect 7267 6218 8067 6248
rect 5533 6216 8067 6218
rect 5533 6160 5538 6216
rect 5594 6160 8067 6216
rect 5533 6158 8067 6160
rect 5533 6155 5599 6158
rect 7267 6128 8067 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 0 5538 800 5568
rect 1301 5538 1367 5541
rect 0 5536 1367 5538
rect 0 5480 1306 5536
rect 1362 5480 1367 5536
rect 0 5478 1367 5480
rect 0 5448 800 5478
rect 1301 5475 1367 5478
rect 6361 5538 6427 5541
rect 7267 5538 8067 5568
rect 6361 5536 8067 5538
rect 6361 5480 6366 5536
rect 6422 5480 8067 5536
rect 6361 5478 8067 5480
rect 6361 5475 6427 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 7267 5448 8067 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 1209 4858 1275 4861
rect 0 4856 1275 4858
rect 0 4800 1214 4856
rect 1270 4800 1275 4856
rect 0 4798 1275 4800
rect 0 4768 800 4798
rect 1209 4795 1275 4798
rect 6177 4858 6243 4861
rect 7267 4858 8067 4888
rect 6177 4856 8067 4858
rect 6177 4800 6182 4856
rect 6238 4800 8067 4856
rect 6177 4798 8067 4800
rect 6177 4795 6243 4798
rect 7267 4768 8067 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4178 800 4208
rect 3233 4178 3299 4181
rect 0 4176 3299 4178
rect 0 4120 3238 4176
rect 3294 4120 3299 4176
rect 0 4118 3299 4120
rect 0 4088 800 4118
rect 3233 4115 3299 4118
rect 5257 4178 5323 4181
rect 7267 4178 8067 4208
rect 5257 4176 8067 4178
rect 5257 4120 5262 4176
rect 5318 4120 8067 4176
rect 5257 4118 8067 4120
rect 5257 4115 5323 4118
rect 7267 4088 8067 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 841 3634 907 3637
rect 798 3632 907 3634
rect 798 3576 846 3632
rect 902 3576 907 3632
rect 798 3571 907 3576
rect 798 3528 858 3571
rect 0 3438 858 3528
rect 6177 3498 6243 3501
rect 7267 3498 8067 3528
rect 6177 3496 8067 3498
rect 6177 3440 6182 3496
rect 6238 3440 8067 3496
rect 6177 3438 8067 3440
rect 0 3408 800 3438
rect 6177 3435 6243 3438
rect 7267 3408 8067 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 5165 2818 5231 2821
rect 7267 2818 8067 2848
rect 5165 2816 8067 2818
rect 5165 2760 5170 2816
rect 5226 2760 8067 2816
rect 5165 2758 8067 2760
rect 5165 2755 5231 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 7267 2728 8067 2758
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 7104 4528 7664
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 7648 5188 7664
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _27_
timestamp 0
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _28_
timestamp 0
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _29_
timestamp 0
transform -1 0 3680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _30_
timestamp 0
transform -1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _31_
timestamp 0
transform -1 0 2024 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _32_
timestamp 0
transform 1 0 1472 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _33_
timestamp 0
transform 1 0 4508 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _34_
timestamp 0
transform -1 0 4784 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _35_
timestamp 0
transform -1 0 5704 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _36_
timestamp 0
transform 1 0 2668 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _37_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _38_
timestamp 0
transform 1 0 3864 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _39_
timestamp 0
transform 1 0 2760 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _40_
timestamp 0
transform -1 0 4324 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _41_
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _42_
timestamp 0
transform -1 0 4968 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _43_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _44_
timestamp 0
transform -1 0 2668 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _45_
timestamp 0
transform -1 0 3864 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _46_
timestamp 0
transform -1 0 3404 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _47_
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _48_
timestamp 0
transform -1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _49_
timestamp 0
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _50_
timestamp 0
transform -1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _51_
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _52_
timestamp 0
transform -1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _53_
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _54_
timestamp 0
transform 1 0 1840 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _55_
timestamp 0
transform 1 0 4784 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _56_
timestamp 0
transform 1 0 1840 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _57_
timestamp 0
transform 1 0 4324 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _58_
timestamp 0
transform -1 0 3404 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _59_
timestamp 0
transform 1 0 4416 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _60_
timestamp 0
transform 1 0 1840 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _61_
timestamp 0
transform 1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 0
transform -1 0 3680 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 0
transform -1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 0
transform -1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 0
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 3220 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_42
timestamp 0
transform 1 0 4968 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 0
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_55
timestamp 0
transform 1 0 6164 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 0
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 0
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_40
timestamp 0
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_16
timestamp 0
transform 1 0 2576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 0
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_38
timestamp 0
transform 1 0 4600 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_50
timestamp 0
transform 1 0 5704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 6256 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 6164 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform 1 0 2024 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform -1 0 4416 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform 1 0 5888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 6624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform -1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform 1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform 1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 0
transform 1 0 5336 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform -1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform 1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 0
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 0
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 0
transform -1 0 3680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 0
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 0
transform -1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_10
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_11
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_12
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_13
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_14
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 6900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_15
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_16
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_17
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_18
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_19
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_22
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_23
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_24
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_25
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_26
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_27
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_28
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_29
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_30
timestamp 0
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_31
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
<< labels >>
rlabel metal1 s 4002 7616 4002 7616 4 VGND
rlabel metal1 s 4002 7072 4002 7072 4 VPWR
rlabel metal2 s 3542 3298 3542 3298 4 _00_
rlabel metal1 s 6578 3162 6578 3162 4 _01_
rlabel metal1 s 3128 5338 3128 5338 4 _02_
rlabel metal1 s 4462 3366 4462 3366 4 _03_
rlabel metal1 s 3128 2618 3128 2618 4 _04_
rlabel metal1 s 6394 2618 6394 2618 4 _05_
rlabel metal2 s 2806 5848 2806 5848 4 _06_
rlabel metal2 s 6486 5202 6486 5202 4 _07_
rlabel metal1 s 2162 3400 2162 3400 4 _08_
rlabel metal2 s 2070 6120 2070 6120 4 _09_
rlabel metal1 s 4738 3162 4738 3162 4 _10_
rlabel metal2 s 3082 3502 3082 3502 4 _11_
rlabel metal1 s 4462 3978 4462 3978 4 _12_
rlabel metal2 s 2162 6494 2162 6494 4 _13_
rlabel metal2 s 4738 6494 4738 6494 4 _14_
rlabel metal2 s 6486 6528 6486 6528 4 _15_
rlabel metal2 s 2346 6647 2346 6647 4 _16_
rlabel metal2 s 3910 4318 3910 4318 4 _17_
rlabel metal1 s 1518 6664 1518 6664 4 _18_
rlabel metal1 s 1978 6426 1978 6426 4 _19_
rlabel metal1 s 4968 6902 4968 6902 4 _20_
rlabel metal1 s 4784 5542 4784 5542 4 _21_
rlabel metal1 s 4462 4794 4462 4794 4 _22_
rlabel metal2 s 3726 3230 3726 3230 4 _23_
rlabel metal1 s 4370 3060 4370 3060 4 _24_
rlabel metal2 s 2622 6324 2622 6324 4 _25_
rlabel metal1 s 3404 4250 3404 4250 4 _26_
rlabel metal2 s 3266 4675 3266 4675 4 clk
rlabel metal1 s 4186 4998 4186 4998 4 clknet_0_clk
rlabel metal1 s 4876 2618 4876 2618 4 clknet_1_0__leaf_clk
rlabel metal2 s 1886 5984 1886 5984 4 clknet_1_1__leaf_clk
rlabel metal1 s 3082 7412 3082 7412 4 eth_data_in[0]
rlabel metal2 s 4554 1588 4554 1588 4 eth_data_in[1]
rlabel metal1 s 1794 7412 1794 7412 4 eth_data_in[2]
rlabel metal3 s 958 4828 958 4828 4 eth_data_in[3]
rlabel metal3 s 1464 8908 1464 8908 4 eth_data_in[4]
rlabel metal1 s 1886 5202 1886 5202 4 eth_data_in[5]
rlabel metal3 s 1004 8228 1004 8228 4 eth_data_in[6]
rlabel metal2 s 5842 7123 5842 7123 4 eth_data_in[7]
rlabel metal1 s 6394 7412 6394 7412 4 eth_valid_in
rlabel metal1 s 4462 5712 4462 5712 4 net1
rlabel metal1 s 3358 2448 3358 2448 4 net10
rlabel metal1 s 1702 5236 1702 5236 4 net11
rlabel metal2 s 6118 3196 6118 3196 4 net12
rlabel metal1 s 5934 2448 5934 2448 4 net13
rlabel metal2 s 1702 3774 1702 3774 4 net14
rlabel metal1 s 5704 5338 5704 5338 4 net15
rlabel metal1 s 2714 7412 2714 7412 4 net16
rlabel metal1 s 4600 2346 4600 2346 4 net17
rlabel metal1 s 2553 7174 2553 7174 4 net18
rlabel metal1 s 5290 6222 5290 6222 4 net19
rlabel metal1 s 4324 2958 4324 2958 4 net2
rlabel metal1 s 1564 5678 1564 5678 4 net20
rlabel metal2 s 6578 4522 6578 4522 4 net21
rlabel metal1 s 5520 4590 5520 4590 4 net22
rlabel metal1 s 4738 2992 4738 2992 4 net23
rlabel metal1 s 2852 4114 2852 4114 4 net24
rlabel metal2 s 2530 6596 2530 6596 4 net25
rlabel metal1 s 2898 6732 2898 6732 4 net26
rlabel metal1 s 6762 6290 6762 6290 4 net27
rlabel metal1 s 3634 4624 3634 4624 4 net28
rlabel metal2 s 1610 7038 1610 7038 4 net3
rlabel metal1 s 1794 6188 1794 6188 4 net4
rlabel metal1 s 2024 5338 2024 5338 4 net5
rlabel metal1 s 1748 5338 1748 5338 4 net6
rlabel metal1 s 2208 7242 2208 7242 4 net7
rlabel metal1 s 1656 6834 1656 6834 4 net8
rlabel metal2 s 5014 7004 5014 7004 4 net9
rlabel metal1 s 1426 5338 1426 5338 4 phy_data_out[0]
rlabel metal3 s 5198 2805 5198 2805 4 phy_data_out[1]
rlabel metal1 s 6164 2618 6164 2618 4 phy_data_out[2]
rlabel metal3 s 0 3408 800 3528 4 phy_data_out[3]
port 16 nsew
rlabel metal2 s 6118 7021 6118 7021 4 phy_data_out[4]
rlabel metal2 s 2622 8476 2622 8476 4 phy_data_out[5]
rlabel metal1 s 5244 4454 5244 4454 4 phy_data_out[6]
rlabel metal1 s 3404 7514 3404 7514 4 phy_data_out[7]
rlabel metal1 s 3680 6630 3680 6630 4 phy_data_out[8]
rlabel metal1 s 1380 5882 1380 5882 4 phy_data_out[9]
rlabel metal2 s 6394 4607 6394 4607 4 phy_valid_out
rlabel metal2 s 6210 4981 6210 4981 4 rst
rlabel metal1 s 4186 4590 4186 4590 4 u_pcs.rd_pos
flabel metal4 s 4868 2128 5188 7664 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4208 2128 4528 7664 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 4088 800 4208 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal2 s 3882 9411 3938 10211 0 FreeSans 280 90 0 0 eth_data_in[0]
port 4 nsew
flabel metal2 s 4526 0 4582 800 0 FreeSans 280 90 0 0 eth_data_in[1]
port 5 nsew
flabel metal2 s 1950 9411 2006 10211 0 FreeSans 280 90 0 0 eth_data_in[2]
port 6 nsew
flabel metal3 s 0 4768 800 4888 0 FreeSans 600 0 0 0 eth_data_in[3]
port 7 nsew
flabel metal3 s 0 8848 800 8968 0 FreeSans 600 0 0 0 eth_data_in[4]
port 8 nsew
flabel metal3 s 0 7488 800 7608 0 FreeSans 600 0 0 0 eth_data_in[5]
port 9 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 eth_data_in[6]
port 10 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 eth_data_in[7]
port 11 nsew
flabel metal2 s 4526 9411 4582 10211 0 FreeSans 280 90 0 0 eth_valid_in
port 12 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 phy_data_out[0]
port 13 nsew
flabel metal3 s 7267 2728 8067 2848 0 FreeSans 600 0 0 0 phy_data_out[1]
port 14 nsew
flabel metal3 s 7267 3408 8067 3528 0 FreeSans 600 0 0 0 phy_data_out[2]
port 15 nsew
flabel metal3 s 400 3468 400 3468 0 FreeSans 600 0 0 0 phy_data_out[3]
flabel metal3 s 7267 6808 8067 6928 0 FreeSans 600 0 0 0 phy_data_out[4]
port 17 nsew
flabel metal2 s 2594 9411 2650 10211 0 FreeSans 280 90 0 0 phy_data_out[5]
port 18 nsew
flabel metal3 s 7267 4088 8067 4208 0 FreeSans 600 0 0 0 phy_data_out[6]
port 19 nsew
flabel metal2 s 3238 9411 3294 10211 0 FreeSans 280 90 0 0 phy_data_out[7]
port 20 nsew
flabel metal3 s 7267 6128 8067 6248 0 FreeSans 600 0 0 0 phy_data_out[8]
port 21 nsew
flabel metal3 s 0 6128 800 6248 0 FreeSans 600 0 0 0 phy_data_out[9]
port 22 nsew
flabel metal3 s 7267 5448 8067 5568 0 FreeSans 600 0 0 0 phy_valid_out
port 23 nsew
flabel metal3 s 7267 4768 8067 4888 0 FreeSans 600 0 0 0 rst
port 24 nsew
<< properties >>
string FIXED_BBOX 0 0 8067 10211
<< end >>
