magic
tech sky130A
magscale 1 2
timestamp 1770939744
<< checkpaint >>
rect -3932 -3932 23236 25380
<< viali >>
rect 8585 18921 8619 18955
rect 9229 18921 9263 18955
rect 11161 18921 11195 18955
rect 11897 18921 11931 18955
rect 8769 18717 8803 18751
rect 9413 18717 9447 18751
rect 11345 18717 11379 18751
rect 11713 18717 11747 18751
rect 11345 14569 11379 14603
rect 1501 14501 1535 14535
rect 1685 14365 1719 14399
rect 5825 14365 5859 14399
rect 9965 14365 9999 14399
rect 14933 14365 14967 14399
rect 15577 14365 15611 14399
rect 16129 14365 16163 14399
rect 17509 14365 17543 14399
rect 10232 14297 10266 14331
rect 6469 14229 6503 14263
rect 14841 14229 14875 14263
rect 17693 14229 17727 14263
rect 1593 14025 1627 14059
rect 4813 14025 4847 14059
rect 6475 14025 6509 14059
rect 6561 14025 6595 14059
rect 6837 14025 6871 14059
rect 8769 14025 8803 14059
rect 9781 14025 9815 14059
rect 11529 14025 11563 14059
rect 14749 14025 14783 14059
rect 16221 14025 16255 14059
rect 17693 14025 17727 14059
rect 5948 13957 5982 13991
rect 9689 13957 9723 13991
rect 1409 13889 1443 13923
rect 6377 13889 6411 13923
rect 6653 13889 6687 13923
rect 6745 13889 6779 13923
rect 7656 13889 7690 13923
rect 9413 13889 9447 13923
rect 9597 13889 9631 13923
rect 9965 13889 9999 13923
rect 10333 13889 10367 13923
rect 12642 13889 12676 13923
rect 12909 13889 12943 13923
rect 13369 13889 13403 13923
rect 13636 13889 13670 13923
rect 14841 13889 14875 13923
rect 15097 13889 15131 13923
rect 17509 13889 17543 13923
rect 6193 13821 6227 13855
rect 7389 13821 7423 13855
rect 10149 13753 10183 13787
rect 8861 13685 8895 13719
rect 9873 13685 9907 13719
rect 6837 13481 6871 13515
rect 10149 13481 10183 13515
rect 10333 13481 10367 13515
rect 13645 13481 13679 13515
rect 13829 13481 13863 13515
rect 14749 13481 14783 13515
rect 8953 13413 8987 13447
rect 9873 13413 9907 13447
rect 6745 13345 6779 13379
rect 6929 13345 6963 13379
rect 11713 13345 11747 13379
rect 1685 13277 1719 13311
rect 7021 13277 7055 13311
rect 9137 13277 9171 13311
rect 9229 13277 9263 13311
rect 9597 13277 9631 13311
rect 9873 13277 9907 13311
rect 14473 13277 14507 13311
rect 14565 13277 14599 13311
rect 14841 13277 14875 13311
rect 15025 13277 15059 13311
rect 17141 13277 17175 13311
rect 17509 13277 17543 13311
rect 10517 13209 10551 13243
rect 13461 13209 13495 13243
rect 14749 13209 14783 13243
rect 14933 13209 14967 13243
rect 1501 13141 1535 13175
rect 9321 13141 9355 13175
rect 9505 13141 9539 13175
rect 10317 13141 10351 13175
rect 12265 13141 12299 13175
rect 13671 13141 13705 13175
rect 17325 13141 17359 13175
rect 17693 13141 17727 13175
rect 6745 12937 6779 12971
rect 7113 12937 7147 12971
rect 8125 12937 8159 12971
rect 9413 12937 9447 12971
rect 9505 12937 9539 12971
rect 9689 12937 9723 12971
rect 13001 12937 13035 12971
rect 13185 12937 13219 12971
rect 6377 12869 6411 12903
rect 6577 12869 6611 12903
rect 6929 12869 6963 12903
rect 7573 12869 7607 12903
rect 10885 12869 10919 12903
rect 11621 12869 11655 12903
rect 12909 12869 12943 12903
rect 15853 12869 15887 12903
rect 16221 12869 16255 12903
rect 1685 12801 1719 12835
rect 6837 12801 6871 12835
rect 7051 12801 7085 12835
rect 7941 12801 7975 12835
rect 8033 12801 8067 12835
rect 8217 12801 8251 12835
rect 9321 12801 9355 12835
rect 10793 12801 10827 12835
rect 11069 12801 11103 12835
rect 11713 12801 11747 12835
rect 12817 12801 12851 12835
rect 15761 12801 15795 12835
rect 16037 12801 16071 12835
rect 16313 12801 16347 12835
rect 16957 12801 16991 12835
rect 7205 12733 7239 12767
rect 7389 12733 7423 12767
rect 7665 12733 7699 12767
rect 7757 12733 7791 12767
rect 7849 12733 7883 12767
rect 9689 12733 9723 12767
rect 13185 12733 13219 12767
rect 17509 12733 17543 12767
rect 11069 12665 11103 12699
rect 1501 12597 1535 12631
rect 6561 12597 6595 12631
rect 16037 12597 16071 12631
rect 7389 12393 7423 12427
rect 9229 12393 9263 12427
rect 14381 12393 14415 12427
rect 17601 12393 17635 12427
rect 6285 12325 6319 12359
rect 13185 12325 13219 12359
rect 6009 12257 6043 12291
rect 7297 12257 7331 12291
rect 11529 12257 11563 12291
rect 13277 12257 13311 12291
rect 14105 12257 14139 12291
rect 4537 12189 4571 12223
rect 5457 12189 5491 12223
rect 5549 12189 5583 12223
rect 5825 12189 5859 12223
rect 6193 12189 6227 12223
rect 6469 12189 6503 12223
rect 7481 12189 7515 12223
rect 7573 12189 7607 12223
rect 11437 12189 11471 12223
rect 11621 12189 11655 12223
rect 11897 12189 11931 12223
rect 12081 12189 12115 12223
rect 12909 12189 12943 12223
rect 14381 12189 14415 12223
rect 14565 12189 14599 12223
rect 14841 12189 14875 12223
rect 15025 12189 15059 12223
rect 15117 12189 15151 12223
rect 15301 12189 15335 12223
rect 16221 12189 16255 12223
rect 6653 12121 6687 12155
rect 9045 12121 9079 12155
rect 11805 12121 11839 12155
rect 13001 12121 13035 12155
rect 16466 12121 16500 12155
rect 4445 12053 4479 12087
rect 6561 12053 6595 12087
rect 6837 12053 6871 12087
rect 9245 12053 9279 12087
rect 9413 12053 9447 12087
rect 11989 12053 12023 12087
rect 13093 12053 13127 12087
rect 14657 12053 14691 12087
rect 15301 12053 15335 12087
rect 4997 11849 5031 11883
rect 6561 11849 6595 11883
rect 6929 11849 6963 11883
rect 9321 11849 9355 11883
rect 9505 11849 9539 11883
rect 10609 11849 10643 11883
rect 13001 11849 13035 11883
rect 5549 11781 5583 11815
rect 6745 11781 6779 11815
rect 8401 11781 8435 11815
rect 1685 11713 1719 11747
rect 3884 11713 3918 11747
rect 5181 11713 5215 11747
rect 5365 11713 5399 11747
rect 6653 11713 6687 11747
rect 8309 11713 8343 11747
rect 8493 11713 8527 11747
rect 8769 11713 8803 11747
rect 8953 11713 8987 11747
rect 9137 11713 9171 11747
rect 9229 11713 9263 11747
rect 9781 11713 9815 11747
rect 10333 11713 10367 11747
rect 10517 11713 10551 11747
rect 11621 11713 11655 11747
rect 11713 11713 11747 11747
rect 11989 11713 12023 11747
rect 12357 11713 12391 11747
rect 12817 11713 12851 11747
rect 14749 11713 14783 11747
rect 15301 11713 15335 11747
rect 15485 11713 15519 11747
rect 15853 11713 15887 11747
rect 16221 11713 16255 11747
rect 16865 11713 16899 11747
rect 3617 11645 3651 11679
rect 9505 11645 9539 11679
rect 9965 11645 9999 11679
rect 16497 11645 16531 11679
rect 17141 11645 17175 11679
rect 6377 11577 6411 11611
rect 10793 11577 10827 11611
rect 16313 11577 16347 11611
rect 17049 11577 17083 11611
rect 1501 11509 1535 11543
rect 8585 11509 8619 11543
rect 9597 11509 9631 11543
rect 11989 11509 12023 11543
rect 14933 11509 14967 11543
rect 16405 11509 16439 11543
rect 16681 11509 16715 11543
rect 4169 11305 4203 11339
rect 7021 11305 7055 11339
rect 11253 11305 11287 11339
rect 12679 11305 12713 11339
rect 15531 11305 15565 11339
rect 15761 11305 15795 11339
rect 17785 11305 17819 11339
rect 5457 11237 5491 11271
rect 10241 11237 10275 11271
rect 12357 11237 12391 11271
rect 15669 11237 15703 11271
rect 12817 11169 12851 11203
rect 14565 11169 14599 11203
rect 14749 11169 14783 11203
rect 14841 11169 14875 11203
rect 4445 11101 4479 11135
rect 4537 11101 4571 11135
rect 4629 11101 4663 11135
rect 4813 11101 4847 11135
rect 4905 11101 4939 11135
rect 5089 11101 5123 11135
rect 5365 11101 5399 11135
rect 5733 11101 5767 11135
rect 6837 11101 6871 11135
rect 9045 11101 9079 11135
rect 9137 11101 9171 11135
rect 9321 11101 9355 11135
rect 9689 11101 9723 11135
rect 9781 11101 9815 11135
rect 9965 11101 9999 11135
rect 10241 11101 10275 11135
rect 11253 11101 11287 11135
rect 11345 11101 11379 11135
rect 12081 11101 12115 11135
rect 12357 11101 12391 11135
rect 12541 11101 12575 11135
rect 13001 11101 13035 11135
rect 14933 11101 14967 11135
rect 15025 11101 15059 11135
rect 15393 11101 15427 11135
rect 15853 11101 15887 11135
rect 16405 11101 16439 11135
rect 16672 11101 16706 11135
rect 4997 11033 5031 11067
rect 6929 11033 6963 11067
rect 7113 11033 7147 11067
rect 10149 11033 10183 11067
rect 11529 11033 11563 11067
rect 12265 11033 12299 11067
rect 5549 10965 5583 10999
rect 5641 10965 5675 10999
rect 13001 10965 13035 10999
rect 5733 10761 5767 10795
rect 6745 10761 6779 10795
rect 14657 10761 14691 10795
rect 14749 10761 14783 10795
rect 1685 10625 1719 10659
rect 3157 10625 3191 10659
rect 5549 10625 5583 10659
rect 5641 10625 5675 10659
rect 6837 10625 6871 10659
rect 6929 10625 6963 10659
rect 10977 10625 11011 10659
rect 12633 10625 12667 10659
rect 14473 10625 14507 10659
rect 14565 10625 14599 10659
rect 17509 10625 17543 10659
rect 5917 10557 5951 10591
rect 6561 10557 6595 10591
rect 14841 10557 14875 10591
rect 5641 10489 5675 10523
rect 1501 10421 1535 10455
rect 2973 10421 3007 10455
rect 6837 10421 6871 10455
rect 10793 10421 10827 10455
rect 13921 10421 13955 10455
rect 17693 10421 17727 10455
rect 3249 10217 3283 10251
rect 5181 10217 5215 10251
rect 8953 10217 8987 10251
rect 11897 10217 11931 10251
rect 17601 10217 17635 10251
rect 13461 10149 13495 10183
rect 3801 10081 3835 10115
rect 5273 10081 5307 10115
rect 6193 10081 6227 10115
rect 7389 10081 7423 10115
rect 10333 10081 10367 10115
rect 13093 10081 13127 10115
rect 16221 10081 16255 10115
rect 1593 10013 1627 10047
rect 1777 10013 1811 10047
rect 1869 10013 1903 10047
rect 5917 10013 5951 10047
rect 6101 10013 6135 10047
rect 6561 10013 6595 10047
rect 7021 10013 7055 10047
rect 7481 10013 7515 10047
rect 7665 10013 7699 10047
rect 7757 10013 7791 10047
rect 7849 10013 7883 10047
rect 8309 10013 8343 10047
rect 8401 10013 8435 10047
rect 10425 10013 10459 10047
rect 10609 10013 10643 10047
rect 10701 10013 10735 10047
rect 10977 10013 11011 10047
rect 11161 10013 11195 10047
rect 11437 10013 11471 10047
rect 11621 10013 11655 10047
rect 11805 10013 11839 10047
rect 11989 10013 12023 10047
rect 12725 10013 12759 10047
rect 12817 10013 12851 10047
rect 13185 10013 13219 10047
rect 13461 10013 13495 10047
rect 13829 10013 13863 10047
rect 15025 10013 15059 10047
rect 15209 10013 15243 10047
rect 16477 10013 16511 10047
rect 1685 9945 1719 9979
rect 2114 9945 2148 9979
rect 4046 9945 4080 9979
rect 6285 9945 6319 9979
rect 6377 9945 6411 9979
rect 8125 9945 8159 9979
rect 10066 9945 10100 9979
rect 11345 9945 11379 9979
rect 6009 9877 6043 9911
rect 7113 9877 7147 9911
rect 7205 9877 7239 9911
rect 7389 9877 7423 9911
rect 12909 9877 12943 9911
rect 13093 9877 13127 9911
rect 13277 9877 13311 9911
rect 13737 9877 13771 9911
rect 15117 9877 15151 9911
rect 3249 9673 3283 9707
rect 3893 9673 3927 9707
rect 5733 9673 5767 9707
rect 5825 9673 5859 9707
rect 8401 9673 8435 9707
rect 13093 9673 13127 9707
rect 13277 9673 13311 9707
rect 13369 9673 13403 9707
rect 14565 9673 14599 9707
rect 1869 9605 1903 9639
rect 2053 9605 2087 9639
rect 2513 9605 2547 9639
rect 12173 9605 12207 9639
rect 14717 9605 14751 9639
rect 14933 9605 14967 9639
rect 1777 9537 1811 9571
rect 2151 9537 2185 9571
rect 3617 9537 3651 9571
rect 4077 9537 4111 9571
rect 5641 9537 5675 9571
rect 6009 9537 6043 9571
rect 8125 9537 8159 9571
rect 8217 9537 8251 9571
rect 8401 9537 8435 9571
rect 9689 9537 9723 9571
rect 9965 9537 9999 9571
rect 10333 9537 10367 9571
rect 10517 9537 10551 9571
rect 10885 9537 10919 9571
rect 11161 9537 11195 9571
rect 11345 9537 11379 9571
rect 12449 9537 12483 9571
rect 12633 9537 12667 9571
rect 12909 9537 12943 9571
rect 13185 9537 13219 9571
rect 14197 9537 14231 9571
rect 14381 9537 14415 9571
rect 14473 9537 14507 9571
rect 15117 9537 15151 9571
rect 15761 9537 15795 9571
rect 16129 9537 16163 9571
rect 16221 9537 16255 9571
rect 17509 9537 17543 9571
rect 3065 9469 3099 9503
rect 3433 9469 3467 9503
rect 3525 9469 3559 9503
rect 3709 9469 3743 9503
rect 4169 9469 4203 9503
rect 4261 9469 4295 9503
rect 9597 9469 9631 9503
rect 12173 9469 12207 9503
rect 12725 9469 12759 9503
rect 13553 9469 13587 9503
rect 2053 9401 2087 9435
rect 2329 9401 2363 9435
rect 6837 9401 6871 9435
rect 11069 9401 11103 9435
rect 12357 9401 12391 9435
rect 12817 9401 12851 9435
rect 14289 9401 14323 9435
rect 17693 9401 17727 9435
rect 5917 9333 5951 9367
rect 13277 9333 13311 9367
rect 14749 9333 14783 9367
rect 15117 9333 15151 9367
rect 6377 9129 6411 9163
rect 12909 9129 12943 9163
rect 15209 9129 15243 9163
rect 17325 9129 17359 9163
rect 9505 9061 9539 9095
rect 5733 8993 5767 9027
rect 8309 8993 8343 9027
rect 8493 8993 8527 9027
rect 12633 8993 12667 9027
rect 12725 8993 12759 9027
rect 15945 8993 15979 9027
rect 5641 8925 5675 8959
rect 5825 8925 5859 8959
rect 5917 8925 5951 8959
rect 8401 8925 8435 8959
rect 8585 8925 8619 8959
rect 9505 8925 9539 8959
rect 9597 8925 9631 8959
rect 10425 8925 10459 8959
rect 10701 8925 10735 8959
rect 12431 8925 12465 8959
rect 12547 8925 12581 8959
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 15025 8925 15059 8959
rect 16201 8925 16235 8959
rect 17509 8925 17543 8959
rect 6193 8857 6227 8891
rect 6409 8857 6443 8891
rect 9781 8857 9815 8891
rect 10609 8857 10643 8891
rect 6101 8789 6135 8823
rect 6561 8789 6595 8823
rect 8125 8789 8159 8823
rect 10885 8789 10919 8823
rect 17693 8789 17727 8823
rect 7481 8585 7515 8619
rect 11161 8585 11195 8619
rect 7665 8517 7699 8551
rect 11805 8517 11839 8551
rect 1869 8449 1903 8483
rect 2237 8449 2271 8483
rect 7389 8449 7423 8483
rect 7757 8449 7791 8483
rect 9045 8449 9079 8483
rect 11069 8449 11103 8483
rect 11621 8449 11655 8483
rect 14105 8449 14139 8483
rect 14289 8449 14323 8483
rect 14657 8449 14691 8483
rect 14749 8449 14783 8483
rect 15025 8449 15059 8483
rect 17509 8449 17543 8483
rect 8033 8381 8067 8415
rect 2053 8313 2087 8347
rect 7665 8313 7699 8347
rect 7849 8313 7883 8347
rect 10333 8313 10367 8347
rect 14841 8313 14875 8347
rect 17693 8313 17727 8347
rect 1685 8245 1719 8279
rect 7757 8245 7791 8279
rect 11989 8245 12023 8279
rect 3157 8041 3191 8075
rect 5457 8041 5491 8075
rect 9045 8041 9079 8075
rect 11253 8041 11287 8075
rect 12633 8041 12667 8075
rect 13001 8041 13035 8075
rect 15025 8041 15059 8075
rect 11069 7973 11103 8007
rect 14749 7973 14783 8007
rect 16589 7973 16623 8007
rect 3617 7905 3651 7939
rect 6837 7905 6871 7939
rect 7205 7905 7239 7939
rect 10149 7905 10183 7939
rect 11345 7905 11379 7939
rect 11437 7905 11471 7939
rect 14841 7905 14875 7939
rect 17417 7905 17451 7939
rect 1685 7837 1719 7871
rect 1777 7837 1811 7871
rect 3433 7837 3467 7871
rect 3801 7837 3835 7871
rect 4169 7837 4203 7871
rect 4721 7837 4755 7871
rect 5089 7837 5123 7871
rect 6570 7837 6604 7871
rect 7472 7837 7506 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 9597 7837 9631 7871
rect 9873 7837 9907 7871
rect 9965 7837 9999 7871
rect 10425 7837 10459 7871
rect 10701 7837 10735 7871
rect 12173 7837 12207 7871
rect 12357 7837 12391 7871
rect 14473 7837 14507 7871
rect 15117 7837 15151 7871
rect 15209 7837 15243 7871
rect 15465 7837 15499 7871
rect 2044 7769 2078 7803
rect 4997 7769 5031 7803
rect 11069 7769 11103 7803
rect 12817 7769 12851 7803
rect 14749 7769 14783 7803
rect 14841 7769 14875 7803
rect 1501 7701 1535 7735
rect 3249 7701 3283 7735
rect 8585 7701 8619 7735
rect 10701 7701 10735 7735
rect 12449 7701 12483 7735
rect 13017 7701 13051 7735
rect 13185 7701 13219 7735
rect 14565 7701 14599 7735
rect 16773 7701 16807 7735
rect 1501 7497 1535 7531
rect 2329 7497 2363 7531
rect 5549 7497 5583 7531
rect 5825 7497 5859 7531
rect 7941 7497 7975 7531
rect 15485 7497 15519 7531
rect 15761 7497 15795 7531
rect 7573 7429 7607 7463
rect 7789 7429 7823 7463
rect 10149 7429 10183 7463
rect 12265 7429 12299 7463
rect 1409 7361 1443 7395
rect 1777 7361 1811 7395
rect 2145 7361 2179 7395
rect 2237 7361 2271 7395
rect 2421 7361 2455 7395
rect 3433 7361 3467 7395
rect 3525 7361 3559 7395
rect 3617 7361 3651 7395
rect 4169 7361 4203 7395
rect 4436 7361 4470 7395
rect 5733 7361 5767 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 10333 7361 10367 7395
rect 10517 7361 10551 7395
rect 10609 7361 10643 7395
rect 11805 7361 11839 7395
rect 11989 7361 12023 7395
rect 14013 7361 14047 7395
rect 14105 7361 14139 7395
rect 14361 7361 14395 7395
rect 15853 7361 15887 7395
rect 1593 7293 1627 7327
rect 3157 7293 3191 7327
rect 3249 7293 3283 7327
rect 3709 7293 3743 7327
rect 1777 7225 1811 7259
rect 2513 7225 2547 7259
rect 1961 7157 1995 7191
rect 7757 7157 7791 7191
rect 10609 7157 10643 7191
rect 11529 7157 11563 7191
rect 11805 7157 11839 7191
rect 4537 6953 4571 6987
rect 10149 6953 10183 6987
rect 11805 6885 11839 6919
rect 12081 6885 12115 6919
rect 3985 6817 4019 6851
rect 9689 6817 9723 6851
rect 1869 6749 1903 6783
rect 2421 6749 2455 6783
rect 2513 6749 2547 6783
rect 3801 6749 3835 6783
rect 4169 6749 4203 6783
rect 4353 6749 4387 6783
rect 4537 6749 4571 6783
rect 4629 6749 4663 6783
rect 4813 6749 4847 6783
rect 9597 6749 9631 6783
rect 9781 6749 9815 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 10609 6749 10643 6783
rect 10793 6749 10827 6783
rect 11713 6749 11747 6783
rect 11805 6749 11839 6783
rect 12357 6749 12391 6783
rect 12541 6749 12575 6783
rect 12817 6749 12851 6783
rect 4721 6681 4755 6715
rect 6653 6681 6687 6715
rect 11529 6681 11563 6715
rect 2605 6613 2639 6647
rect 3893 6613 3927 6647
rect 4077 6613 4111 6647
rect 10793 6613 10827 6647
rect 12265 6613 12299 6647
rect 1593 6409 1627 6443
rect 3233 6409 3267 6443
rect 9413 6409 9447 6443
rect 3433 6341 3467 6375
rect 8125 6341 8159 6375
rect 2706 6273 2740 6307
rect 8309 6273 8343 6307
rect 8585 6273 8619 6307
rect 8769 6273 8803 6307
rect 9045 6273 9079 6307
rect 9137 6273 9171 6307
rect 9321 6273 9355 6307
rect 9689 6273 9723 6307
rect 9781 6273 9815 6307
rect 10517 6273 10551 6307
rect 10885 6273 10919 6307
rect 11069 6273 11103 6307
rect 2973 6205 3007 6239
rect 9505 6205 9539 6239
rect 10425 6205 10459 6239
rect 9689 6137 9723 6171
rect 3065 6069 3099 6103
rect 3249 6069 3283 6103
rect 6837 6069 6871 6103
rect 10701 6069 10735 6103
rect 10885 6069 10919 6103
rect 2145 5865 2179 5899
rect 2605 5865 2639 5899
rect 13645 5865 13679 5899
rect 7757 5797 7791 5831
rect 11897 5797 11931 5831
rect 2973 5729 3007 5763
rect 3065 5729 3099 5763
rect 3249 5729 3283 5763
rect 11713 5729 11747 5763
rect 1869 5661 1903 5695
rect 1961 5661 1995 5695
rect 2329 5661 2363 5695
rect 2532 5661 2566 5695
rect 2697 5661 2731 5695
rect 3157 5661 3191 5695
rect 4169 5661 4203 5695
rect 4261 5661 4295 5695
rect 4353 5661 4387 5695
rect 4629 5661 4663 5695
rect 6101 5661 6135 5695
rect 6285 5661 6319 5695
rect 6377 5661 6411 5695
rect 8401 5661 8435 5695
rect 8769 5661 8803 5695
rect 9137 5661 9171 5695
rect 9413 5661 9447 5695
rect 10802 5661 10836 5695
rect 11069 5661 11103 5695
rect 11529 5661 11563 5695
rect 11621 5661 11655 5695
rect 11897 5661 11931 5695
rect 11989 5661 12023 5695
rect 12173 5661 12207 5695
rect 12265 5661 12299 5695
rect 2145 5593 2179 5627
rect 4537 5593 4571 5627
rect 4874 5593 4908 5627
rect 6193 5593 6227 5627
rect 6622 5593 6656 5627
rect 7849 5593 7883 5627
rect 9229 5593 9263 5627
rect 12510 5593 12544 5627
rect 2421 5525 2455 5559
rect 2789 5525 2823 5559
rect 3985 5525 4019 5559
rect 6009 5525 6043 5559
rect 8677 5525 8711 5559
rect 9597 5525 9631 5559
rect 9689 5525 9723 5559
rect 12081 5525 12115 5559
rect 3617 5321 3651 5355
rect 4169 5321 4203 5355
rect 6745 5321 6779 5355
rect 7021 5321 7055 5355
rect 8401 5321 8435 5355
rect 8677 5321 8711 5355
rect 12265 5321 12299 5355
rect 4997 5253 5031 5287
rect 7205 5253 7239 5287
rect 7573 5253 7607 5287
rect 7757 5253 7791 5287
rect 3525 5185 3559 5219
rect 3893 5185 3927 5219
rect 4077 5185 4111 5219
rect 4261 5185 4295 5219
rect 4629 5185 4663 5219
rect 4813 5185 4847 5219
rect 6653 5185 6687 5219
rect 6837 5185 6871 5219
rect 6929 5185 6963 5219
rect 7297 5185 7331 5219
rect 7665 5185 7699 5219
rect 7941 5185 7975 5219
rect 8125 5185 8159 5219
rect 8217 5185 8251 5219
rect 8309 5185 8343 5219
rect 8585 5185 8619 5219
rect 12265 5185 12299 5219
rect 12449 5185 12483 5219
rect 3709 5117 3743 5151
rect 4353 5117 4387 5151
rect 4537 5117 4571 5151
rect 4721 5117 4755 5151
rect 5549 5117 5583 5151
rect 7481 5117 7515 5151
rect 9229 5117 9263 5151
rect 3893 5049 3927 5083
rect 7297 5049 7331 5083
rect 8309 5049 8343 5083
rect 7205 4981 7239 5015
rect 13369 4777 13403 4811
rect 12817 4709 12851 4743
rect 9229 4641 9263 4675
rect 12449 4641 12483 4675
rect 7389 4573 7423 4607
rect 7645 4573 7679 4607
rect 9137 4573 9171 4607
rect 9321 4573 9355 4607
rect 9413 4573 9447 4607
rect 13093 4573 13127 4607
rect 13185 4573 13219 4607
rect 17785 4573 17819 4607
rect 12633 4505 12667 4539
rect 12817 4505 12851 4539
rect 8769 4437 8803 4471
rect 8953 4437 8987 4471
rect 13001 4437 13035 4471
rect 17601 4437 17635 4471
rect 4261 4233 4295 4267
rect 5917 4233 5951 4267
rect 6561 4233 6595 4267
rect 6929 4233 6963 4267
rect 10057 4233 10091 4267
rect 10149 4233 10183 4267
rect 11713 4233 11747 4267
rect 11989 4233 12023 4267
rect 8125 4165 8159 4199
rect 11805 4165 11839 4199
rect 12808 4165 12842 4199
rect 4169 4097 4203 4131
rect 4537 4097 4571 4131
rect 4721 4097 4755 4131
rect 4905 4097 4939 4131
rect 5641 4097 5675 4131
rect 6009 4097 6043 4131
rect 6101 4097 6135 4131
rect 6653 4097 6687 4131
rect 6745 4097 6779 4131
rect 7113 4097 7147 4131
rect 7205 4097 7239 4131
rect 7389 4097 7423 4131
rect 7849 4097 7883 4131
rect 7941 4097 7975 4131
rect 9965 4097 9999 4131
rect 11897 4097 11931 4131
rect 12173 4097 12207 4131
rect 12357 4097 12391 4131
rect 12541 4097 12575 4131
rect 4353 4029 4387 4063
rect 4997 4029 5031 4063
rect 5733 4029 5767 4063
rect 6377 4029 6411 4063
rect 10333 4029 10367 4063
rect 11069 4029 11103 4063
rect 11529 4029 11563 4063
rect 14565 4029 14599 4063
rect 7297 3961 7331 3995
rect 10057 3961 10091 3995
rect 13921 3961 13955 3995
rect 4537 3893 4571 3927
rect 4813 3893 4847 3927
rect 5825 3893 5859 3927
rect 6653 3893 6687 3927
rect 8125 3893 8159 3927
rect 10425 3893 10459 3927
rect 11805 3893 11839 3927
rect 14013 3893 14047 3927
rect 7941 3689 7975 3723
rect 9045 3689 9079 3723
rect 10609 3689 10643 3723
rect 12541 3689 12575 3723
rect 12817 3689 12851 3723
rect 5641 3621 5675 3655
rect 9505 3621 9539 3655
rect 4445 3485 4479 3519
rect 4629 3485 4663 3519
rect 5365 3485 5399 3519
rect 5641 3485 5675 3519
rect 5733 3485 5767 3519
rect 7757 3485 7791 3519
rect 8125 3485 8159 3519
rect 8217 3485 8251 3519
rect 8769 3485 8803 3519
rect 9137 3485 9171 3519
rect 9505 3485 9539 3519
rect 9781 3485 9815 3519
rect 10241 3485 10275 3519
rect 10701 3485 10735 3519
rect 11161 3485 11195 3519
rect 11529 3485 11563 3519
rect 11897 3485 11931 3519
rect 12357 3485 12391 3519
rect 12449 3485 12483 3519
rect 12633 3485 12667 3519
rect 12909 3485 12943 3519
rect 5978 3417 6012 3451
rect 12081 3417 12115 3451
rect 4537 3349 4571 3383
rect 5457 3349 5491 3383
rect 7113 3349 7147 3383
rect 7205 3349 7239 3383
rect 8585 3349 8619 3383
rect 9689 3349 9723 3383
rect 10149 3349 10183 3383
rect 12179 3349 12213 3383
rect 12265 3349 12299 3383
rect 6469 3145 6503 3179
rect 9137 3145 9171 3179
rect 10609 3145 10643 3179
rect 11621 3145 11655 3179
rect 4160 3077 4194 3111
rect 9496 3077 9530 3111
rect 10961 3077 10995 3111
rect 11161 3077 11195 3111
rect 3893 3009 3927 3043
rect 6561 3009 6595 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 7481 3009 7515 3043
rect 8217 3009 8251 3043
rect 11529 3009 11563 3043
rect 11713 3009 11747 3043
rect 12918 3009 12952 3043
rect 13185 3009 13219 3043
rect 8585 2941 8619 2975
rect 9229 2941 9263 2975
rect 10793 2873 10827 2907
rect 5273 2805 5307 2839
rect 8125 2805 8159 2839
rect 10977 2805 11011 2839
rect 11805 2805 11839 2839
rect 13553 2601 13587 2635
rect 8769 2533 8803 2567
rect 12817 2533 12851 2567
rect 7389 2465 7423 2499
rect 12633 2465 12667 2499
rect 5549 2397 5583 2431
rect 5917 2397 5951 2431
rect 6929 2397 6963 2431
rect 7297 2397 7331 2431
rect 7656 2397 7690 2431
rect 9137 2397 9171 2431
rect 9781 2397 9815 2431
rect 10425 2397 10459 2431
rect 11069 2397 11103 2431
rect 11897 2397 11931 2431
rect 11989 2397 12023 2431
rect 13001 2397 13035 2431
rect 13369 2397 13403 2431
rect 13461 2397 13495 2431
rect 5733 2261 5767 2295
rect 6101 2261 6135 2295
rect 6745 2261 6779 2295
rect 7113 2261 7147 2295
rect 9321 2261 9355 2295
rect 9965 2261 9999 2295
rect 10609 2261 10643 2295
rect 11253 2261 11287 2295
rect 11713 2261 11747 2295
rect 13185 2261 13219 2295
<< metal1 >>
rect 1104 19066 18124 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 18124 19066
rect 1104 18992 18124 19014
rect 8570 18912 8576 18964
rect 8628 18912 8634 18964
rect 9214 18912 9220 18964
rect 9272 18912 9278 18964
rect 10870 18912 10876 18964
rect 10928 18952 10934 18964
rect 11149 18955 11207 18961
rect 11149 18952 11161 18955
rect 10928 18924 11161 18952
rect 10928 18912 10934 18924
rect 11149 18921 11161 18924
rect 11195 18921 11207 18955
rect 11149 18915 11207 18921
rect 11882 18912 11888 18964
rect 11940 18912 11946 18964
rect 8754 18708 8760 18760
rect 8812 18708 8818 18760
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18748 9459 18751
rect 9582 18748 9588 18760
rect 9447 18720 9588 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 11330 18708 11336 18760
rect 11388 18708 11394 18760
rect 11698 18708 11704 18760
rect 11756 18708 11762 18760
rect 1104 18522 18124 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 18124 18522
rect 1104 18448 18124 18470
rect 1104 17978 18124 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 18124 17978
rect 1104 17904 18124 17926
rect 1104 17434 18124 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 18124 17434
rect 1104 17360 18124 17382
rect 1104 16890 18124 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 18124 16890
rect 1104 16816 18124 16838
rect 1104 16346 18124 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 18124 16346
rect 1104 16272 18124 16294
rect 1104 15802 18124 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 18124 15802
rect 1104 15728 18124 15750
rect 1104 15258 18124 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 18124 15258
rect 1104 15184 18124 15206
rect 1104 14714 18124 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 18124 14714
rect 1104 14640 18124 14662
rect 11330 14560 11336 14612
rect 11388 14560 11394 14612
rect 842 14492 848 14544
rect 900 14532 906 14544
rect 1489 14535 1547 14541
rect 1489 14532 1501 14535
rect 900 14504 1501 14532
rect 900 14492 906 14504
rect 1489 14501 1501 14504
rect 1535 14501 1547 14535
rect 1489 14495 1547 14501
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 4798 14396 4804 14408
rect 1719 14368 4804 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 4798 14356 4804 14368
rect 4856 14396 4862 14408
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 4856 14368 5825 14396
rect 4856 14356 4862 14368
rect 5813 14365 5825 14368
rect 5859 14396 5871 14399
rect 6270 14396 6276 14408
rect 5859 14368 6276 14396
rect 5859 14365 5871 14368
rect 5813 14359 5871 14365
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 9953 14399 10011 14405
rect 9953 14365 9965 14399
rect 9999 14396 10011 14399
rect 12894 14396 12900 14408
rect 9999 14368 12900 14396
rect 9999 14365 10011 14368
rect 9953 14359 10011 14365
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 14921 14399 14979 14405
rect 14921 14365 14933 14399
rect 14967 14396 14979 14399
rect 15565 14399 15623 14405
rect 15565 14396 15577 14399
rect 14967 14368 15577 14396
rect 14967 14365 14979 14368
rect 14921 14359 14979 14365
rect 15565 14365 15577 14368
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 16114 14356 16120 14408
rect 16172 14396 16178 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 16172 14368 17509 14396
rect 16172 14356 16178 14368
rect 17497 14365 17509 14368
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 10226 14337 10232 14340
rect 10220 14291 10232 14337
rect 10226 14288 10232 14291
rect 10284 14288 10290 14340
rect 6457 14263 6515 14269
rect 6457 14229 6469 14263
rect 6503 14260 6515 14263
rect 6730 14260 6736 14272
rect 6503 14232 6736 14260
rect 6503 14229 6515 14232
rect 6457 14223 6515 14229
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 14550 14220 14556 14272
rect 14608 14260 14614 14272
rect 14829 14263 14887 14269
rect 14829 14260 14841 14263
rect 14608 14232 14841 14260
rect 14608 14220 14614 14232
rect 14829 14229 14841 14232
rect 14875 14229 14887 14263
rect 14829 14223 14887 14229
rect 17678 14220 17684 14272
rect 17736 14220 17742 14272
rect 1104 14170 18124 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 18124 14170
rect 1104 14096 18124 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 2130 14056 2136 14068
rect 1627 14028 2136 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 2130 14016 2136 14028
rect 2188 14016 2194 14068
rect 4798 14016 4804 14068
rect 4856 14016 4862 14068
rect 6463 14059 6521 14065
rect 6463 14056 6475 14059
rect 6196 14028 6475 14056
rect 5936 13991 5994 13997
rect 5936 13957 5948 13991
rect 5982 13988 5994 13991
rect 6196 13988 6224 14028
rect 6463 14025 6475 14028
rect 6509 14025 6521 14059
rect 6463 14019 6521 14025
rect 6549 14059 6607 14065
rect 6549 14025 6561 14059
rect 6595 14056 6607 14059
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6595 14028 6837 14056
rect 6595 14025 6607 14028
rect 6549 14019 6607 14025
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 6825 14019 6883 14025
rect 8754 14016 8760 14068
rect 8812 14016 8818 14068
rect 8938 14016 8944 14068
rect 8996 14056 9002 14068
rect 9769 14059 9827 14065
rect 9769 14056 9781 14059
rect 8996 14028 9781 14056
rect 8996 14016 9002 14028
rect 9769 14025 9781 14028
rect 9815 14056 9827 14059
rect 11330 14056 11336 14068
rect 9815 14028 11336 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11698 14056 11704 14068
rect 11563 14028 11704 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 7098 13988 7104 14000
rect 5982 13960 6224 13988
rect 6656 13960 7104 13988
rect 5982 13957 5994 13960
rect 5936 13951 5994 13957
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 6362 13880 6368 13932
rect 6420 13880 6426 13932
rect 6656 13929 6684 13960
rect 7098 13948 7104 13960
rect 7156 13948 7162 14000
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 6730 13880 6736 13932
rect 6788 13880 6794 13932
rect 7644 13923 7702 13929
rect 7644 13889 7656 13923
rect 7690 13920 7702 13923
rect 8110 13920 8116 13932
rect 7690 13892 8116 13920
rect 7690 13889 7702 13892
rect 7644 13883 7702 13889
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 8772 13920 8800 14016
rect 9677 13991 9735 13997
rect 9677 13988 9689 13991
rect 9416 13960 9689 13988
rect 9122 13920 9128 13932
rect 8772 13892 9128 13920
rect 9122 13880 9128 13892
rect 9180 13920 9186 13932
rect 9416 13929 9444 13960
rect 9677 13957 9689 13960
rect 9723 13957 9735 13991
rect 11532 13988 11560 14019
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 14792 14028 15332 14056
rect 14792 14016 14798 14028
rect 15194 13988 15200 14000
rect 9677 13951 9735 13957
rect 9968 13960 11560 13988
rect 13372 13960 15200 13988
rect 9968 13932 9996 13960
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 9180 13892 9413 13920
rect 9180 13880 9186 13892
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 9582 13880 9588 13932
rect 9640 13880 9646 13932
rect 9950 13880 9956 13932
rect 10008 13880 10014 13932
rect 10318 13880 10324 13932
rect 10376 13880 10382 13932
rect 12618 13880 12624 13932
rect 12676 13929 12682 13932
rect 12676 13883 12688 13929
rect 12676 13880 12682 13883
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 13372 13929 13400 13960
rect 13357 13923 13415 13929
rect 13357 13920 13369 13923
rect 12952 13892 13369 13920
rect 12952 13880 12958 13892
rect 13357 13889 13369 13892
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13624 13923 13682 13929
rect 13624 13889 13636 13923
rect 13670 13920 13682 13923
rect 13906 13920 13912 13932
rect 13670 13892 13912 13920
rect 13670 13889 13682 13892
rect 13624 13883 13682 13889
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 14844 13929 14872 13960
rect 15194 13948 15200 13960
rect 15252 13948 15258 14000
rect 15304 13988 15332 14028
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 16114 14056 16120 14068
rect 15528 14028 16120 14056
rect 15528 14016 15534 14028
rect 16114 14016 16120 14028
rect 16172 14056 16178 14068
rect 16209 14059 16267 14065
rect 16209 14056 16221 14059
rect 16172 14028 16221 14056
rect 16172 14016 16178 14028
rect 16209 14025 16221 14028
rect 16255 14025 16267 14059
rect 16209 14019 16267 14025
rect 17678 14016 17684 14068
rect 17736 14016 17742 14068
rect 15304 13960 16574 13988
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 14918 13880 14924 13932
rect 14976 13920 14982 13932
rect 15085 13923 15143 13929
rect 15085 13920 15097 13923
rect 14976 13892 15097 13920
rect 14976 13880 14982 13892
rect 15085 13889 15097 13892
rect 15131 13889 15143 13923
rect 16546 13920 16574 13960
rect 17497 13923 17555 13929
rect 17497 13920 17509 13923
rect 16546 13892 17509 13920
rect 15085 13883 15143 13889
rect 17497 13889 17509 13892
rect 17543 13889 17555 13923
rect 17497 13883 17555 13889
rect 6181 13855 6239 13861
rect 6181 13821 6193 13855
rect 6227 13852 6239 13855
rect 6914 13852 6920 13864
rect 6227 13824 6920 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 6914 13812 6920 13824
rect 6972 13852 6978 13864
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 6972 13824 7389 13852
rect 6972 13812 6978 13824
rect 7377 13821 7389 13824
rect 7423 13821 7435 13855
rect 7377 13815 7435 13821
rect 9306 13744 9312 13796
rect 9364 13784 9370 13796
rect 10137 13787 10195 13793
rect 10137 13784 10149 13787
rect 9364 13756 10149 13784
rect 9364 13744 9370 13756
rect 10137 13753 10149 13756
rect 10183 13784 10195 13787
rect 11146 13784 11152 13796
rect 10183 13756 11152 13784
rect 10183 13753 10195 13756
rect 10137 13747 10195 13753
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 8846 13676 8852 13728
rect 8904 13676 8910 13728
rect 9858 13676 9864 13728
rect 9916 13676 9922 13728
rect 1104 13626 18124 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 18124 13626
rect 1104 13552 18124 13574
rect 6362 13472 6368 13524
rect 6420 13512 6426 13524
rect 6825 13515 6883 13521
rect 6825 13512 6837 13515
rect 6420 13484 6837 13512
rect 6420 13472 6426 13484
rect 6825 13481 6837 13484
rect 6871 13481 6883 13515
rect 6825 13475 6883 13481
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 10226 13512 10232 13524
rect 10183 13484 10232 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 10321 13515 10379 13521
rect 10321 13481 10333 13515
rect 10367 13512 10379 13515
rect 10367 13484 12940 13512
rect 10367 13481 10379 13484
rect 10321 13475 10379 13481
rect 8938 13404 8944 13456
rect 8996 13404 9002 13456
rect 9861 13447 9919 13453
rect 9861 13413 9873 13447
rect 9907 13444 9919 13447
rect 12066 13444 12072 13456
rect 9907 13416 12072 13444
rect 9907 13413 9919 13416
rect 9861 13407 9919 13413
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 6546 13336 6552 13388
rect 6604 13376 6610 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 6604 13348 6745 13376
rect 6604 13336 6610 13348
rect 6733 13345 6745 13348
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7466 13376 7472 13388
rect 6963 13348 7472 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 11698 13336 11704 13388
rect 11756 13336 11762 13388
rect 12912 13376 12940 13484
rect 12986 13472 12992 13524
rect 13044 13512 13050 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 13044 13484 13645 13512
rect 13044 13472 13050 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 13633 13475 13691 13481
rect 13817 13515 13875 13521
rect 13817 13481 13829 13515
rect 13863 13512 13875 13515
rect 13906 13512 13912 13524
rect 13863 13484 13912 13512
rect 13863 13481 13875 13484
rect 13817 13475 13875 13481
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 14737 13515 14795 13521
rect 14737 13481 14749 13515
rect 14783 13512 14795 13515
rect 14918 13512 14924 13524
rect 14783 13484 14924 13512
rect 14783 13481 14795 13484
rect 14737 13475 14795 13481
rect 14918 13472 14924 13484
rect 14976 13472 14982 13524
rect 13630 13376 13636 13388
rect 12912 13348 13636 13376
rect 13630 13336 13636 13348
rect 13688 13376 13694 13388
rect 13688 13348 15056 13376
rect 13688 13336 13694 13348
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 4614 13308 4620 13320
rect 1719 13280 4620 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 7064 13280 9076 13308
rect 7064 13268 7070 13280
rect 9048 13240 9076 13280
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9490 13308 9496 13320
rect 9272 13280 9496 13308
rect 9272 13268 9278 13280
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 9585 13311 9643 13317
rect 9585 13277 9597 13311
rect 9631 13277 9643 13311
rect 9585 13271 9643 13277
rect 9600 13240 9628 13271
rect 9858 13268 9864 13320
rect 9916 13268 9922 13320
rect 11882 13308 11888 13320
rect 10428 13280 11888 13308
rect 10428 13240 10456 13280
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 9048 13212 10456 13240
rect 10502 13200 10508 13252
rect 10560 13200 10566 13252
rect 13446 13200 13452 13252
rect 13504 13240 13510 13252
rect 14476 13240 14504 13271
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 14826 13268 14832 13320
rect 14884 13268 14890 13320
rect 15028 13317 15056 13348
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13308 15071 13311
rect 15838 13308 15844 13320
rect 15059 13280 15844 13308
rect 15059 13277 15071 13280
rect 15013 13271 15071 13277
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 17126 13268 17132 13320
rect 17184 13268 17190 13320
rect 17494 13268 17500 13320
rect 17552 13268 17558 13320
rect 13504 13212 14504 13240
rect 14737 13243 14795 13249
rect 13504 13200 13510 13212
rect 14737 13209 14749 13243
rect 14783 13240 14795 13243
rect 14921 13243 14979 13249
rect 14921 13240 14933 13243
rect 14783 13212 14933 13240
rect 14783 13209 14795 13212
rect 14737 13203 14795 13209
rect 14921 13209 14933 13212
rect 14967 13209 14979 13243
rect 14921 13203 14979 13209
rect 842 13132 848 13184
rect 900 13172 906 13184
rect 1489 13175 1547 13181
rect 1489 13172 1501 13175
rect 900 13144 1501 13172
rect 900 13132 906 13144
rect 1489 13141 1501 13144
rect 1535 13141 1547 13175
rect 1489 13135 1547 13141
rect 9306 13132 9312 13184
rect 9364 13132 9370 13184
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 9456 13144 9505 13172
rect 9456 13132 9462 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9493 13135 9551 13141
rect 10305 13175 10363 13181
rect 10305 13141 10317 13175
rect 10351 13172 10363 13175
rect 10594 13172 10600 13184
rect 10351 13144 10600 13172
rect 10351 13141 10363 13144
rect 10305 13135 10363 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 12253 13175 12311 13181
rect 12253 13172 12265 13175
rect 11756 13144 12265 13172
rect 11756 13132 11762 13144
rect 12253 13141 12265 13144
rect 12299 13141 12311 13175
rect 12253 13135 12311 13141
rect 13659 13175 13717 13181
rect 13659 13141 13671 13175
rect 13705 13172 13717 13175
rect 14366 13172 14372 13184
rect 13705 13144 14372 13172
rect 13705 13141 13717 13144
rect 13659 13135 13717 13141
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 17310 13132 17316 13184
rect 17368 13132 17374 13184
rect 17678 13132 17684 13184
rect 17736 13132 17742 13184
rect 1104 13082 18124 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 18124 13082
rect 1104 13008 18124 13030
rect 6733 12971 6791 12977
rect 6733 12937 6745 12971
rect 6779 12937 6791 12971
rect 6733 12931 6791 12937
rect 6362 12860 6368 12912
rect 6420 12860 6426 12912
rect 6565 12903 6623 12909
rect 6565 12900 6577 12903
rect 6472 12872 6577 12900
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 5534 12832 5540 12844
rect 1719 12804 5540 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 5534 12792 5540 12804
rect 5592 12832 5598 12844
rect 6472 12832 6500 12872
rect 6565 12869 6577 12872
rect 6611 12869 6623 12903
rect 6565 12863 6623 12869
rect 5592 12804 6500 12832
rect 6748 12832 6776 12931
rect 7098 12928 7104 12980
rect 7156 12928 7162 12980
rect 8110 12928 8116 12980
rect 8168 12928 8174 12980
rect 9398 12928 9404 12980
rect 9456 12928 9462 12980
rect 9490 12928 9496 12980
rect 9548 12928 9554 12980
rect 9677 12971 9735 12977
rect 9677 12937 9689 12971
rect 9723 12937 9735 12971
rect 9677 12931 9735 12937
rect 12989 12971 13047 12977
rect 12989 12937 13001 12971
rect 13035 12937 13047 12971
rect 12989 12931 13047 12937
rect 13173 12971 13231 12977
rect 13173 12937 13185 12971
rect 13219 12968 13231 12971
rect 13446 12968 13452 12980
rect 13219 12940 13452 12968
rect 13219 12937 13231 12940
rect 13173 12931 13231 12937
rect 6917 12903 6975 12909
rect 6917 12869 6929 12903
rect 6963 12900 6975 12903
rect 7561 12903 7619 12909
rect 7561 12900 7573 12903
rect 6963 12872 7573 12900
rect 6963 12869 6975 12872
rect 6917 12863 6975 12869
rect 7561 12869 7573 12872
rect 7607 12900 7619 12903
rect 9508 12900 9536 12928
rect 7607 12872 9536 12900
rect 9692 12900 9720 12931
rect 10502 12900 10508 12912
rect 9692 12872 10508 12900
rect 7607 12869 7619 12872
rect 7561 12863 7619 12869
rect 10502 12860 10508 12872
rect 10560 12900 10566 12912
rect 10873 12903 10931 12909
rect 10560 12872 10824 12900
rect 10560 12860 10566 12872
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6748 12804 6837 12832
rect 5592 12792 5598 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 7039 12835 7097 12841
rect 7039 12801 7051 12835
rect 7085 12832 7097 12835
rect 7929 12835 7987 12841
rect 7085 12804 7420 12832
rect 7085 12801 7097 12804
rect 7039 12795 7097 12801
rect 7392 12773 7420 12804
rect 7929 12801 7941 12835
rect 7975 12832 7987 12835
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7975 12804 8033 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 8021 12801 8033 12804
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 8202 12792 8208 12844
rect 8260 12792 8266 12844
rect 9306 12792 9312 12844
rect 9364 12792 9370 12844
rect 10796 12841 10824 12872
rect 10873 12869 10885 12903
rect 10919 12900 10931 12903
rect 11514 12900 11520 12912
rect 10919 12872 11520 12900
rect 10919 12869 10931 12872
rect 10873 12863 10931 12869
rect 11514 12860 11520 12872
rect 11572 12900 11578 12912
rect 11609 12903 11667 12909
rect 11609 12900 11621 12903
rect 11572 12872 11621 12900
rect 11572 12860 11578 12872
rect 11609 12869 11621 12872
rect 11655 12869 11667 12903
rect 11609 12863 11667 12869
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 12897 12903 12955 12909
rect 12897 12900 12909 12903
rect 12124 12872 12909 12900
rect 12124 12860 12130 12872
rect 12897 12869 12909 12872
rect 12943 12869 12955 12903
rect 13004 12900 13032 12931
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 13262 12900 13268 12912
rect 13004 12872 13268 12900
rect 12897 12863 12955 12869
rect 13262 12860 13268 12872
rect 13320 12860 13326 12912
rect 15841 12903 15899 12909
rect 15841 12869 15853 12903
rect 15887 12900 15899 12903
rect 16209 12903 16267 12909
rect 16209 12900 16221 12903
rect 15887 12872 16221 12900
rect 15887 12869 15899 12872
rect 15841 12863 15899 12869
rect 16209 12869 16221 12872
rect 16255 12869 16267 12903
rect 16209 12863 16267 12869
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 11054 12792 11060 12844
rect 11112 12792 11118 12844
rect 11698 12792 11704 12844
rect 11756 12792 11762 12844
rect 12802 12792 12808 12844
rect 12860 12792 12866 12844
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 14884 12804 15761 12832
rect 14884 12792 14890 12804
rect 15749 12801 15761 12804
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15988 12804 16037 12832
rect 15988 12792 15994 12804
rect 16025 12801 16037 12804
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16347 12804 16957 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 7377 12767 7435 12773
rect 7377 12733 7389 12767
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 7208 12640 7236 12727
rect 7392 12696 7420 12727
rect 7650 12724 7656 12776
rect 7708 12724 7714 12776
rect 7742 12724 7748 12776
rect 7800 12724 7806 12776
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 8846 12764 8852 12776
rect 7883 12736 8852 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 8846 12724 8852 12736
rect 8904 12724 8910 12776
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 10226 12764 10232 12776
rect 9723 12736 10232 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 9692 12696 9720 12727
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12764 13231 12767
rect 14734 12764 14740 12776
rect 13219 12736 14740 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 17494 12724 17500 12776
rect 17552 12724 17558 12776
rect 7392 12668 9720 12696
rect 11057 12699 11115 12705
rect 11057 12665 11069 12699
rect 11103 12696 11115 12699
rect 12618 12696 12624 12708
rect 11103 12668 12624 12696
rect 11103 12665 11115 12668
rect 11057 12659 11115 12665
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 1486 12588 1492 12640
rect 1544 12588 1550 12640
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12628 6607 12631
rect 6638 12628 6644 12640
rect 6595 12600 6644 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 7190 12588 7196 12640
rect 7248 12628 7254 12640
rect 7742 12628 7748 12640
rect 7248 12600 7748 12628
rect 7248 12588 7254 12600
rect 7742 12588 7748 12600
rect 7800 12628 7806 12640
rect 10318 12628 10324 12640
rect 7800 12600 10324 12628
rect 7800 12588 7806 12600
rect 10318 12588 10324 12600
rect 10376 12628 10382 12640
rect 13814 12628 13820 12640
rect 10376 12600 13820 12628
rect 10376 12588 10382 12600
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 16022 12588 16028 12640
rect 16080 12588 16086 12640
rect 1104 12538 18124 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 18124 12538
rect 1104 12464 18124 12486
rect 6362 12424 6368 12436
rect 5828 12396 6368 12424
rect 5828 12288 5856 12396
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 7377 12427 7435 12433
rect 7377 12393 7389 12427
rect 7423 12424 7435 12427
rect 8202 12424 8208 12436
rect 7423 12396 8208 12424
rect 7423 12393 7435 12396
rect 7377 12387 7435 12393
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 9030 12384 9036 12436
rect 9088 12424 9094 12436
rect 9217 12427 9275 12433
rect 9217 12424 9229 12427
rect 9088 12396 9229 12424
rect 9088 12384 9094 12396
rect 9217 12393 9229 12396
rect 9263 12393 9275 12427
rect 9217 12387 9275 12393
rect 14366 12384 14372 12436
rect 14424 12384 14430 12436
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 17589 12427 17647 12433
rect 17589 12424 17601 12427
rect 17552 12396 17601 12424
rect 17552 12384 17558 12396
rect 17589 12393 17601 12396
rect 17635 12393 17647 12427
rect 17589 12387 17647 12393
rect 6270 12316 6276 12368
rect 6328 12316 6334 12368
rect 6546 12316 6552 12368
rect 6604 12356 6610 12368
rect 13173 12359 13231 12365
rect 6604 12328 7328 12356
rect 6604 12316 6610 12328
rect 4632 12260 5856 12288
rect 4632 12232 4660 12260
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12220 4583 12223
rect 4614 12220 4620 12232
rect 4571 12192 4620 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 5445 12223 5503 12229
rect 5445 12189 5457 12223
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 5460 12152 5488 12183
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 5828 12229 5856 12260
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12288 6055 12291
rect 7006 12288 7012 12300
rect 6043 12260 7012 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7300 12297 7328 12328
rect 13173 12325 13185 12359
rect 13219 12356 13231 12359
rect 14826 12356 14832 12368
rect 13219 12328 14832 12356
rect 13219 12325 13231 12328
rect 13173 12319 13231 12325
rect 14826 12316 14832 12328
rect 14884 12316 14890 12368
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12288 7343 12291
rect 7742 12288 7748 12300
rect 7331 12260 7748 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 11514 12248 11520 12300
rect 11572 12288 11578 12300
rect 11572 12260 12112 12288
rect 11572 12248 11578 12260
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6270 12220 6276 12232
rect 6227 12192 6276 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 6362 12180 6368 12232
rect 6420 12220 6426 12232
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 6420 12192 6469 12220
rect 6420 12180 6426 12192
rect 6457 12189 6469 12192
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 7466 12180 7472 12232
rect 7524 12180 7530 12232
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12220 7619 12223
rect 8386 12220 8392 12232
rect 7607 12192 8392 12220
rect 7607 12189 7619 12192
rect 7561 12183 7619 12189
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 11422 12180 11428 12232
rect 11480 12180 11486 12232
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12220 11667 12223
rect 11882 12220 11888 12232
rect 11655 12192 11888 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 12084 12229 12112 12260
rect 13262 12248 13268 12300
rect 13320 12248 13326 12300
rect 14093 12291 14151 12297
rect 14093 12257 14105 12291
rect 14139 12288 14151 12291
rect 14458 12288 14464 12300
rect 14139 12260 14464 12288
rect 14139 12257 14151 12260
rect 14093 12251 14151 12257
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 14660 12260 15148 12288
rect 12069 12223 12127 12229
rect 12069 12189 12081 12223
rect 12115 12189 12127 12223
rect 12069 12183 12127 12189
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 12897 12223 12955 12229
rect 12897 12220 12909 12223
rect 12860 12192 12909 12220
rect 12860 12180 12866 12192
rect 12897 12189 12909 12192
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 14366 12180 14372 12232
rect 14424 12180 14430 12232
rect 14550 12180 14556 12232
rect 14608 12180 14614 12232
rect 5626 12152 5632 12164
rect 5460 12124 5632 12152
rect 5626 12112 5632 12124
rect 5684 12152 5690 12164
rect 6641 12155 6699 12161
rect 6641 12152 6653 12155
rect 5684 12124 6653 12152
rect 5684 12112 5690 12124
rect 6641 12121 6653 12124
rect 6687 12121 6699 12155
rect 6641 12115 6699 12121
rect 8938 12112 8944 12164
rect 8996 12152 9002 12164
rect 9033 12155 9091 12161
rect 9033 12152 9045 12155
rect 8996 12124 9045 12152
rect 8996 12112 9002 12124
rect 9033 12121 9045 12124
rect 9079 12152 9091 12155
rect 9582 12152 9588 12164
rect 9079 12124 9588 12152
rect 9079 12121 9091 12124
rect 9033 12115 9091 12121
rect 9582 12112 9588 12124
rect 9640 12112 9646 12164
rect 11793 12155 11851 12161
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 12986 12152 12992 12164
rect 11839 12124 12992 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 4433 12087 4491 12093
rect 4433 12053 4445 12087
rect 4479 12084 4491 12087
rect 4614 12084 4620 12096
rect 4479 12056 4620 12084
rect 4479 12053 4491 12056
rect 4433 12047 4491 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 6546 12084 6552 12096
rect 5500 12056 6552 12084
rect 5500 12044 5506 12056
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 6825 12087 6883 12093
rect 6825 12053 6837 12087
rect 6871 12084 6883 12087
rect 7006 12084 7012 12096
rect 6871 12056 7012 12084
rect 6871 12053 6883 12056
rect 6825 12047 6883 12053
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 8754 12044 8760 12096
rect 8812 12084 8818 12096
rect 9214 12084 9220 12096
rect 9272 12093 9278 12096
rect 9272 12087 9291 12093
rect 8812 12056 9220 12084
rect 8812 12044 8818 12056
rect 9214 12044 9220 12056
rect 9279 12053 9291 12087
rect 9272 12047 9291 12053
rect 9272 12044 9278 12047
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 11422 12084 11428 12096
rect 9456 12056 11428 12084
rect 9456 12044 9462 12056
rect 11422 12044 11428 12056
rect 11480 12044 11486 12096
rect 11606 12044 11612 12096
rect 11664 12084 11670 12096
rect 14660 12093 14688 12260
rect 14826 12180 14832 12232
rect 14884 12180 14890 12232
rect 15120 12229 15148 12260
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15252 12260 16252 12288
rect 15252 12248 15258 12260
rect 16224 12232 16252 12260
rect 15013 12223 15071 12229
rect 15013 12189 15025 12223
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12189 15163 12223
rect 15105 12183 15163 12189
rect 15028 12152 15056 12183
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15344 12192 15976 12220
rect 15344 12180 15350 12192
rect 15470 12152 15476 12164
rect 15028 12124 15476 12152
rect 15470 12112 15476 12124
rect 15528 12112 15534 12164
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11664 12056 11989 12084
rect 11664 12044 11670 12056
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 11977 12047 12035 12053
rect 13081 12087 13139 12093
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 13127 12056 14657 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 14645 12053 14657 12056
rect 14691 12084 14703 12087
rect 14734 12084 14740 12096
rect 14691 12056 14740 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15289 12087 15347 12093
rect 15289 12053 15301 12087
rect 15335 12084 15347 12087
rect 15378 12084 15384 12096
rect 15335 12056 15384 12084
rect 15335 12053 15347 12056
rect 15289 12047 15347 12053
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 15948 12084 15976 12192
rect 16206 12180 16212 12232
rect 16264 12180 16270 12232
rect 16022 12112 16028 12164
rect 16080 12152 16086 12164
rect 16454 12155 16512 12161
rect 16454 12152 16466 12155
rect 16080 12124 16466 12152
rect 16080 12112 16086 12124
rect 16454 12121 16466 12124
rect 16500 12121 16512 12155
rect 16454 12115 16512 12121
rect 17494 12084 17500 12096
rect 15948 12056 17500 12084
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 1104 11994 18124 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 18124 11994
rect 1104 11920 18124 11942
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4764 11852 4997 11880
rect 4764 11840 4770 11852
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 4985 11843 5043 11849
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6328 11852 6561 11880
rect 6328 11840 6334 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 6549 11843 6607 11849
rect 6917 11883 6975 11889
rect 6917 11849 6929 11883
rect 6963 11880 6975 11883
rect 7650 11880 7656 11892
rect 6963 11852 7656 11880
rect 6963 11849 6975 11852
rect 6917 11843 6975 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 8754 11880 8760 11892
rect 8352 11852 8760 11880
rect 8352 11840 8358 11852
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 9309 11883 9367 11889
rect 9309 11880 9321 11883
rect 9272 11852 9321 11880
rect 9272 11840 9278 11852
rect 9309 11849 9321 11852
rect 9355 11849 9367 11883
rect 9309 11843 9367 11849
rect 9490 11840 9496 11892
rect 9548 11840 9554 11892
rect 10594 11840 10600 11892
rect 10652 11840 10658 11892
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 12989 11883 13047 11889
rect 12989 11880 13001 11883
rect 12860 11852 13001 11880
rect 12860 11840 12866 11852
rect 12989 11849 13001 11852
rect 13035 11849 13047 11883
rect 12989 11843 13047 11849
rect 15838 11840 15844 11892
rect 15896 11840 15902 11892
rect 5442 11812 5448 11824
rect 1688 11784 5448 11812
rect 1688 11753 1716 11784
rect 3878 11753 3884 11756
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 3872 11707 3884 11753
rect 3878 11704 3884 11707
rect 3936 11704 3942 11756
rect 5184 11753 5212 11784
rect 5442 11772 5448 11784
rect 5500 11772 5506 11824
rect 5537 11815 5595 11821
rect 5537 11781 5549 11815
rect 5583 11812 5595 11815
rect 5718 11812 5724 11824
rect 5583 11784 5724 11812
rect 5583 11781 5595 11784
rect 5537 11775 5595 11781
rect 5718 11772 5724 11784
rect 5776 11812 5782 11824
rect 6733 11815 6791 11821
rect 6733 11812 6745 11815
rect 5776 11784 6745 11812
rect 5776 11772 5782 11784
rect 6733 11781 6745 11784
rect 6779 11781 6791 11815
rect 6733 11775 6791 11781
rect 8386 11772 8392 11824
rect 8444 11812 8450 11824
rect 8662 11812 8668 11824
rect 8444 11784 8668 11812
rect 8444 11772 8450 11784
rect 8662 11772 8668 11784
rect 8720 11772 8726 11824
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11744 5411 11747
rect 5626 11744 5632 11756
rect 5399 11716 5632 11744
rect 5399 11713 5411 11716
rect 5353 11707 5411 11713
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 6420 11716 6653 11744
rect 6420 11704 6426 11716
rect 6641 11713 6653 11716
rect 6687 11713 6699 11747
rect 6641 11707 6699 11713
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 8202 11744 8208 11756
rect 7064 11716 8208 11744
rect 7064 11704 7070 11716
rect 8202 11704 8208 11716
rect 8260 11744 8266 11756
rect 8772 11753 8800 11840
rect 9398 11812 9404 11824
rect 9140 11784 9404 11812
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 8260 11716 8309 11744
rect 8260 11704 8266 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11744 8539 11747
rect 8757 11747 8815 11753
rect 8527 11716 8616 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 3602 11636 3608 11688
rect 3660 11636 3666 11688
rect 6365 11611 6423 11617
rect 6365 11577 6377 11611
rect 6411 11608 6423 11611
rect 8294 11608 8300 11620
rect 6411 11580 8300 11608
rect 6411 11577 6423 11580
rect 6365 11571 6423 11577
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 842 11500 848 11552
rect 900 11540 906 11552
rect 8588 11549 8616 11716
rect 8757 11713 8769 11747
rect 8803 11713 8815 11747
rect 8757 11707 8815 11713
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11744 8999 11747
rect 9030 11744 9036 11756
rect 8987 11716 9036 11744
rect 8987 11713 8999 11716
rect 8941 11707 8999 11713
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9140 11753 9168 11784
rect 9398 11772 9404 11784
rect 9456 11772 9462 11824
rect 9508 11784 10364 11812
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11713 9183 11747
rect 9125 11707 9183 11713
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9306 11744 9312 11756
rect 9263 11716 9312 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 9508 11744 9536 11784
rect 9416 11716 9536 11744
rect 8662 11568 8668 11620
rect 8720 11608 8726 11620
rect 9416 11608 9444 11716
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9640 11716 9781 11744
rect 9640 11704 9646 11716
rect 9769 11713 9781 11716
rect 9815 11744 9827 11747
rect 10042 11744 10048 11756
rect 9815 11716 10048 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 10336 11753 10364 11784
rect 11422 11772 11428 11824
rect 11480 11812 11486 11824
rect 11480 11784 11744 11812
rect 11480 11772 11486 11784
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11744 10563 11747
rect 11238 11744 11244 11756
rect 10551 11716 11244 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11606 11704 11612 11756
rect 11664 11704 11670 11756
rect 11716 11753 11744 11784
rect 14826 11772 14832 11824
rect 14884 11812 14890 11824
rect 15856 11812 15884 11840
rect 14884 11784 15608 11812
rect 15856 11784 16896 11812
rect 14884 11772 14890 11784
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11974 11704 11980 11756
rect 12032 11704 12038 11756
rect 12342 11704 12348 11756
rect 12400 11704 12406 11756
rect 12802 11704 12808 11756
rect 12860 11704 12866 11756
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11744 14795 11747
rect 14918 11744 14924 11756
rect 14783 11716 14924 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 15286 11704 15292 11756
rect 15344 11704 15350 11756
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15580 11744 15608 11784
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 15580 11716 15853 11744
rect 15841 11713 15853 11716
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 16868 11753 16896 11784
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 16172 11716 16221 11744
rect 16172 11704 16178 11716
rect 16209 11713 16221 11716
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11645 9551 11679
rect 9950 11676 9956 11688
rect 9493 11639 9551 11645
rect 9646 11648 9956 11676
rect 8720 11580 9444 11608
rect 9508 11608 9536 11639
rect 9646 11608 9674 11648
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 16485 11679 16543 11685
rect 16485 11676 16497 11679
rect 15436 11648 16497 11676
rect 15436 11636 15442 11648
rect 16485 11645 16497 11648
rect 16531 11645 16543 11679
rect 16485 11639 16543 11645
rect 17126 11636 17132 11688
rect 17184 11676 17190 11688
rect 17770 11676 17776 11688
rect 17184 11648 17776 11676
rect 17184 11636 17190 11648
rect 17770 11636 17776 11648
rect 17828 11636 17834 11688
rect 9508 11580 9674 11608
rect 8720 11568 8726 11580
rect 10042 11568 10048 11620
rect 10100 11608 10106 11620
rect 10781 11611 10839 11617
rect 10781 11608 10793 11611
rect 10100 11580 10793 11608
rect 10100 11568 10106 11580
rect 10781 11577 10793 11580
rect 10827 11577 10839 11611
rect 10781 11571 10839 11577
rect 14550 11568 14556 11620
rect 14608 11608 14614 11620
rect 16301 11611 16359 11617
rect 16301 11608 16313 11611
rect 14608 11580 16313 11608
rect 14608 11568 14614 11580
rect 16301 11577 16313 11580
rect 16347 11577 16359 11611
rect 17037 11611 17095 11617
rect 17037 11608 17049 11611
rect 16301 11571 16359 11577
rect 16408 11580 17049 11608
rect 1489 11543 1547 11549
rect 1489 11540 1501 11543
rect 900 11512 1501 11540
rect 900 11500 906 11512
rect 1489 11509 1501 11512
rect 1535 11509 1547 11543
rect 1489 11503 1547 11509
rect 8573 11543 8631 11549
rect 8573 11509 8585 11543
rect 8619 11540 8631 11543
rect 9398 11540 9404 11552
rect 8619 11512 9404 11540
rect 8619 11509 8631 11512
rect 8573 11503 8631 11509
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9585 11543 9643 11549
rect 9585 11509 9597 11543
rect 9631 11540 9643 11543
rect 9766 11540 9772 11552
rect 9631 11512 9772 11540
rect 9631 11509 9643 11512
rect 9585 11503 9643 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 11977 11543 12035 11549
rect 11977 11509 11989 11543
rect 12023 11540 12035 11543
rect 12066 11540 12072 11552
rect 12023 11512 12072 11540
rect 12023 11509 12035 11512
rect 11977 11503 12035 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 16408 11549 16436 11580
rect 17037 11577 17049 11580
rect 17083 11577 17095 11611
rect 17037 11571 17095 11577
rect 14921 11543 14979 11549
rect 14921 11540 14933 11543
rect 14884 11512 14933 11540
rect 14884 11500 14890 11512
rect 14921 11509 14933 11512
rect 14967 11509 14979 11543
rect 14921 11503 14979 11509
rect 16393 11543 16451 11549
rect 16393 11509 16405 11543
rect 16439 11509 16451 11543
rect 16393 11503 16451 11509
rect 16666 11500 16672 11552
rect 16724 11500 16730 11552
rect 1104 11450 18124 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 18124 11450
rect 1104 11376 18124 11398
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 4157 11339 4215 11345
rect 4157 11336 4169 11339
rect 3936 11308 4169 11336
rect 3936 11296 3942 11308
rect 4157 11305 4169 11308
rect 4203 11305 4215 11339
rect 4157 11299 4215 11305
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 6454 11336 6460 11348
rect 4764 11308 6460 11336
rect 4764 11296 4770 11308
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 7009 11339 7067 11345
rect 7009 11305 7021 11339
rect 7055 11336 7067 11339
rect 7466 11336 7472 11348
rect 7055 11308 7472 11336
rect 7055 11305 7067 11308
rect 7009 11299 7067 11305
rect 7466 11296 7472 11308
rect 7524 11296 7530 11348
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 12667 11339 12725 11345
rect 12667 11336 12679 11339
rect 11296 11308 12679 11336
rect 11296 11296 11302 11308
rect 12667 11305 12679 11308
rect 12713 11305 12725 11339
rect 12667 11299 12725 11305
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 15519 11339 15577 11345
rect 15519 11336 15531 11339
rect 14608 11308 15531 11336
rect 14608 11296 14614 11308
rect 15519 11305 15531 11308
rect 15565 11305 15577 11339
rect 15519 11299 15577 11305
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11336 15807 11339
rect 15930 11336 15936 11348
rect 15795 11308 15936 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 17770 11296 17776 11348
rect 17828 11296 17834 11348
rect 4614 11228 4620 11280
rect 4672 11268 4678 11280
rect 5445 11271 5503 11277
rect 4672 11240 4844 11268
rect 4672 11228 4678 11240
rect 4632 11200 4660 11228
rect 4448 11172 4660 11200
rect 4816 11200 4844 11240
rect 5445 11237 5457 11271
rect 5491 11237 5503 11271
rect 9674 11268 9680 11280
rect 5445 11231 5503 11237
rect 9232 11240 9680 11268
rect 5460 11200 5488 11231
rect 9232 11212 9260 11240
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 10229 11271 10287 11277
rect 10229 11237 10241 11271
rect 10275 11237 10287 11271
rect 10229 11231 10287 11237
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11268 12403 11271
rect 14366 11268 14372 11280
rect 12391 11240 14372 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 9214 11200 9220 11212
rect 4816 11172 4936 11200
rect 4448 11141 4476 11172
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4522 11092 4528 11144
rect 4580 11092 4586 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 4706 11132 4712 11144
rect 4663 11104 4712 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 4908 11141 4936 11172
rect 5092 11172 5488 11200
rect 9048 11172 9220 11200
rect 5092 11141 5120 11172
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 4816 11064 4844 11095
rect 4985 11067 5043 11073
rect 4985 11064 4997 11067
rect 4816 11036 4997 11064
rect 4985 11033 4997 11036
rect 5031 11033 5043 11067
rect 5368 11064 5396 11095
rect 5718 11092 5724 11144
rect 5776 11092 5782 11144
rect 6546 11092 6552 11144
rect 6604 11132 6610 11144
rect 9048 11141 9076 11172
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 9490 11200 9496 11212
rect 9324 11172 9496 11200
rect 6825 11135 6883 11141
rect 6825 11132 6837 11135
rect 6604 11104 6837 11132
rect 6604 11092 6610 11104
rect 6825 11101 6837 11104
rect 6871 11101 6883 11135
rect 6825 11095 6883 11101
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 9324 11141 9352 11172
rect 9490 11160 9496 11172
rect 9548 11200 9554 11212
rect 10244 11200 10272 11231
rect 14366 11228 14372 11240
rect 14424 11268 14430 11280
rect 15657 11271 15715 11277
rect 15657 11268 15669 11271
rect 14424 11240 15669 11268
rect 14424 11228 14430 11240
rect 15657 11237 15669 11240
rect 15703 11268 15715 11271
rect 16114 11268 16120 11280
rect 15703 11240 16120 11268
rect 15703 11237 15715 11240
rect 15657 11231 15715 11237
rect 16114 11228 16120 11240
rect 16172 11228 16178 11280
rect 12805 11203 12863 11209
rect 9548 11172 10088 11200
rect 10244 11172 12572 11200
rect 9548 11160 9554 11172
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9456 11104 9689 11132
rect 9456 11092 9462 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 6564 11064 6592 11092
rect 5368 11036 6592 11064
rect 4985 11027 5043 11033
rect 6730 11024 6736 11076
rect 6788 11064 6794 11076
rect 6917 11067 6975 11073
rect 6917 11064 6929 11067
rect 6788 11036 6929 11064
rect 6788 11024 6794 11036
rect 6917 11033 6929 11036
rect 6963 11033 6975 11067
rect 6917 11027 6975 11033
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11033 7159 11067
rect 9692 11064 9720 11095
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9824 11104 9965 11132
rect 9824 11092 9830 11104
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 10060 11132 10088 11172
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 10060 11104 10241 11132
rect 9953 11095 10011 11101
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 11146 11092 11152 11144
rect 11204 11132 11210 11144
rect 11241 11135 11299 11141
rect 11241 11132 11253 11135
rect 11204 11104 11253 11132
rect 11204 11092 11210 11104
rect 11241 11101 11253 11104
rect 11287 11101 11299 11135
rect 11241 11095 11299 11101
rect 11330 11092 11336 11144
rect 11388 11092 11394 11144
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11132 12127 11135
rect 12158 11132 12164 11144
rect 12115 11104 12164 11132
rect 12115 11101 12127 11104
rect 12069 11095 12127 11101
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 12544 11141 12572 11172
rect 12805 11169 12817 11203
rect 12851 11200 12863 11203
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 12851 11172 14565 11200
rect 12851 11169 12863 11172
rect 12805 11163 12863 11169
rect 14553 11169 14565 11172
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 14734 11160 14740 11212
rect 14792 11160 14798 11212
rect 14829 11203 14887 11209
rect 14829 11169 14841 11203
rect 14875 11200 14887 11203
rect 15286 11200 15292 11212
rect 14875 11172 15292 11200
rect 14875 11169 14887 11172
rect 14829 11163 14887 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12676 11104 13001 11132
rect 12676 11092 12682 11104
rect 12989 11101 13001 11104
rect 13035 11132 13047 11135
rect 13078 11132 13084 11144
rect 13035 11104 13084 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 14918 11092 14924 11144
rect 14976 11092 14982 11144
rect 15010 11092 15016 11144
rect 15068 11092 15074 11144
rect 15378 11092 15384 11144
rect 15436 11092 15442 11144
rect 15838 11092 15844 11144
rect 15896 11092 15902 11144
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 16666 11141 16672 11144
rect 16393 11135 16451 11141
rect 16393 11132 16405 11135
rect 16264 11104 16405 11132
rect 16264 11092 16270 11104
rect 16393 11101 16405 11104
rect 16439 11101 16451 11135
rect 16660 11132 16672 11141
rect 16627 11104 16672 11132
rect 16393 11095 16451 11101
rect 16660 11095 16672 11104
rect 16666 11092 16672 11095
rect 16724 11092 16730 11144
rect 10137 11067 10195 11073
rect 10137 11064 10149 11067
rect 9692 11036 10149 11064
rect 7101 11027 7159 11033
rect 10137 11033 10149 11036
rect 10183 11033 10195 11067
rect 10137 11027 10195 11033
rect 5534 10956 5540 11008
rect 5592 10956 5598 11008
rect 5629 10999 5687 11005
rect 5629 10965 5641 10999
rect 5675 10996 5687 10999
rect 6822 10996 6828 11008
rect 5675 10968 6828 10996
rect 5675 10965 5687 10968
rect 5629 10959 5687 10965
rect 6822 10956 6828 10968
rect 6880 10996 6886 11008
rect 7116 10996 7144 11027
rect 10686 11024 10692 11076
rect 10744 11064 10750 11076
rect 11517 11067 11575 11073
rect 11517 11064 11529 11067
rect 10744 11036 11529 11064
rect 10744 11024 10750 11036
rect 11517 11033 11529 11036
rect 11563 11064 11575 11067
rect 11974 11064 11980 11076
rect 11563 11036 11980 11064
rect 11563 11033 11575 11036
rect 11517 11027 11575 11033
rect 11974 11024 11980 11036
rect 12032 11064 12038 11076
rect 12253 11067 12311 11073
rect 12253 11064 12265 11067
rect 12032 11036 12265 11064
rect 12032 11024 12038 11036
rect 12253 11033 12265 11036
rect 12299 11033 12311 11067
rect 12253 11027 12311 11033
rect 6880 10968 7144 10996
rect 6880 10956 6886 10968
rect 10410 10956 10416 11008
rect 10468 10996 10474 11008
rect 11330 10996 11336 11008
rect 10468 10968 11336 10996
rect 10468 10956 10474 10968
rect 11330 10956 11336 10968
rect 11388 10996 11394 11008
rect 12360 10996 12388 11092
rect 14936 11064 14964 11092
rect 17126 11064 17132 11076
rect 14936 11036 17132 11064
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 11388 10968 12388 10996
rect 12989 10999 13047 11005
rect 11388 10956 11394 10968
rect 12989 10965 13001 10999
rect 13035 10996 13047 10999
rect 13446 10996 13452 11008
rect 13035 10968 13452 10996
rect 13035 10965 13047 10968
rect 12989 10959 13047 10965
rect 13446 10956 13452 10968
rect 13504 10956 13510 11008
rect 1104 10906 18124 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 18124 10906
rect 1104 10832 18124 10854
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5721 10795 5779 10801
rect 5721 10792 5733 10795
rect 5592 10764 5733 10792
rect 5592 10752 5598 10764
rect 5721 10761 5733 10764
rect 5767 10792 5779 10795
rect 6730 10792 6736 10804
rect 5767 10764 6736 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 14550 10752 14556 10804
rect 14608 10792 14614 10804
rect 14645 10795 14703 10801
rect 14645 10792 14657 10795
rect 14608 10764 14657 10792
rect 14608 10752 14614 10764
rect 14645 10761 14657 10764
rect 14691 10761 14703 10795
rect 14645 10755 14703 10761
rect 14734 10752 14740 10804
rect 14792 10752 14798 10804
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 3050 10656 3056 10668
rect 1719 10628 3056 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 3050 10616 3056 10628
rect 3108 10616 3114 10668
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10656 3203 10659
rect 3510 10656 3516 10668
rect 3191 10628 3516 10656
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 6822 10656 6828 10668
rect 5675 10628 6828 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5552 10588 5580 10619
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7006 10656 7012 10668
rect 6963 10628 7012 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10744 10628 10977 10656
rect 10744 10616 10750 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 12492 10628 12633 10656
rect 12492 10616 12498 10628
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14458 10656 14464 10668
rect 13872 10628 14464 10656
rect 13872 10616 13878 10628
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 14553 10659 14611 10665
rect 14553 10625 14565 10659
rect 14599 10656 14611 10659
rect 15102 10656 15108 10668
rect 14599 10628 15108 10656
rect 14599 10625 14611 10628
rect 14553 10619 14611 10625
rect 15102 10616 15108 10628
rect 15160 10656 15166 10668
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 15160 10628 17509 10656
rect 15160 10616 15166 10628
rect 17497 10625 17509 10628
rect 17543 10656 17555 10659
rect 17586 10656 17592 10668
rect 17543 10628 17592 10656
rect 17543 10625 17555 10628
rect 17497 10619 17555 10625
rect 17586 10616 17592 10628
rect 17644 10616 17650 10668
rect 5718 10588 5724 10600
rect 5552 10560 5724 10588
rect 5718 10548 5724 10560
rect 5776 10548 5782 10600
rect 5902 10548 5908 10600
rect 5960 10548 5966 10600
rect 6546 10548 6552 10600
rect 6604 10548 6610 10600
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 14826 10588 14832 10600
rect 14424 10560 14832 10588
rect 14424 10548 14430 10560
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 4522 10480 4528 10532
rect 4580 10520 4586 10532
rect 5629 10523 5687 10529
rect 5629 10520 5641 10523
rect 4580 10492 5641 10520
rect 4580 10480 4586 10492
rect 5629 10489 5641 10492
rect 5675 10489 5687 10523
rect 5629 10483 5687 10489
rect 842 10412 848 10464
rect 900 10452 906 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 900 10424 1501 10452
rect 900 10412 906 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 1489 10415 1547 10421
rect 2958 10412 2964 10464
rect 3016 10412 3022 10464
rect 6825 10455 6883 10461
rect 6825 10421 6837 10455
rect 6871 10452 6883 10455
rect 8202 10452 8208 10464
rect 6871 10424 8208 10452
rect 6871 10421 6883 10424
rect 6825 10415 6883 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10376 10424 10793 10452
rect 10376 10412 10382 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 12158 10452 12164 10464
rect 11204 10424 12164 10452
rect 11204 10412 11210 10424
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 12768 10424 13921 10452
rect 12768 10412 12774 10424
rect 13909 10421 13921 10424
rect 13955 10452 13967 10455
rect 16206 10452 16212 10464
rect 13955 10424 16212 10452
rect 13955 10421 13967 10424
rect 13909 10415 13967 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 17678 10412 17684 10464
rect 17736 10412 17742 10464
rect 1104 10362 18124 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 18124 10362
rect 1104 10288 18124 10310
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3237 10251 3295 10257
rect 3237 10248 3249 10251
rect 3108 10220 3249 10248
rect 3108 10208 3114 10220
rect 3237 10217 3249 10220
rect 3283 10217 3295 10251
rect 3237 10211 3295 10217
rect 5169 10251 5227 10257
rect 5169 10217 5181 10251
rect 5215 10248 5227 10251
rect 5442 10248 5448 10260
rect 5215 10220 5448 10248
rect 5215 10217 5227 10220
rect 5169 10211 5227 10217
rect 3602 10072 3608 10124
rect 3660 10112 3666 10124
rect 5276 10121 5304 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8812 10220 8953 10248
rect 8812 10208 8818 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 8941 10211 8999 10217
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 11885 10251 11943 10257
rect 11885 10248 11897 10251
rect 11112 10220 11897 10248
rect 11112 10208 11118 10220
rect 11885 10217 11897 10220
rect 11931 10217 11943 10251
rect 11885 10211 11943 10217
rect 12894 10208 12900 10260
rect 12952 10248 12958 10260
rect 14550 10248 14556 10260
rect 12952 10220 14556 10248
rect 12952 10208 12958 10220
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 17586 10208 17592 10260
rect 17644 10208 17650 10260
rect 5902 10140 5908 10192
rect 5960 10180 5966 10192
rect 9122 10180 9128 10192
rect 5960 10152 9128 10180
rect 5960 10140 5966 10152
rect 3789 10115 3847 10121
rect 3789 10112 3801 10115
rect 3660 10084 3801 10112
rect 3660 10072 3666 10084
rect 3789 10081 3801 10084
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10081 5319 10115
rect 5261 10075 5319 10081
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6822 10112 6828 10124
rect 6227 10084 6828 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 7392 10121 7420 10152
rect 9122 10140 9128 10152
rect 9180 10140 9186 10192
rect 12710 10180 12716 10192
rect 12406 10152 12716 10180
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10081 7435 10115
rect 8478 10112 8484 10124
rect 7377 10075 7435 10081
rect 7484 10084 8484 10112
rect 1578 10004 1584 10056
rect 1636 10004 1642 10056
rect 1762 10004 1768 10056
rect 1820 10004 1826 10056
rect 1854 10004 1860 10056
rect 1912 10044 1918 10056
rect 3620 10044 3648 10072
rect 1912 10016 3648 10044
rect 5905 10047 5963 10053
rect 1912 10004 1918 10016
rect 5905 10013 5917 10047
rect 5951 10044 5963 10047
rect 6089 10047 6147 10053
rect 6089 10044 6101 10047
rect 5951 10016 6101 10044
rect 5951 10013 5963 10016
rect 5905 10007 5963 10013
rect 6089 10013 6101 10016
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 7006 10004 7012 10056
rect 7064 10004 7070 10056
rect 7484 10053 7512 10084
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 10321 10115 10379 10121
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 12406 10112 12434 10152
rect 12710 10140 12716 10152
rect 12768 10140 12774 10192
rect 13262 10140 13268 10192
rect 13320 10140 13326 10192
rect 13449 10183 13507 10189
rect 13449 10149 13461 10183
rect 13495 10180 13507 10183
rect 13495 10152 15332 10180
rect 13495 10149 13507 10152
rect 13449 10143 13507 10149
rect 10367 10084 12434 10112
rect 13081 10115 13139 10121
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 13081 10081 13093 10115
rect 13127 10112 13139 10115
rect 13280 10112 13308 10140
rect 13127 10084 13308 10112
rect 13127 10081 13139 10084
rect 13081 10075 13139 10081
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7650 10004 7656 10056
rect 7708 10004 7714 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8294 10044 8300 10056
rect 7883 10016 8300 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 2102 9979 2160 9985
rect 2102 9976 2114 9979
rect 1719 9948 2114 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 2102 9945 2114 9948
rect 2148 9945 2160 9979
rect 2102 9939 2160 9945
rect 3878 9936 3884 9988
rect 3936 9976 3942 9988
rect 4034 9979 4092 9985
rect 4034 9976 4046 9979
rect 3936 9948 4046 9976
rect 3936 9936 3942 9948
rect 4034 9945 4046 9948
rect 4080 9945 4092 9979
rect 4034 9939 4092 9945
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 6273 9979 6331 9985
rect 6273 9976 6285 9979
rect 5684 9948 6285 9976
rect 5684 9936 5690 9948
rect 6273 9945 6285 9948
rect 6319 9945 6331 9979
rect 6273 9939 6331 9945
rect 6365 9979 6423 9985
rect 6365 9945 6377 9979
rect 6411 9976 6423 9979
rect 6730 9976 6736 9988
rect 6411 9948 6736 9976
rect 6411 9945 6423 9948
rect 6365 9939 6423 9945
rect 6730 9936 6736 9948
rect 6788 9976 6794 9988
rect 7760 9976 7788 10007
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10044 8447 10047
rect 8754 10044 8760 10056
rect 8435 10016 8760 10044
rect 8435 10013 8447 10016
rect 8389 10007 8447 10013
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10594 10004 10600 10056
rect 10652 10004 10658 10056
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10796 10016 10977 10044
rect 6788 9948 7236 9976
rect 6788 9936 6794 9948
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 5997 9911 6055 9917
rect 5997 9908 6009 9911
rect 5592 9880 6009 9908
rect 5592 9868 5598 9880
rect 5997 9877 6009 9880
rect 6043 9877 6055 9911
rect 5997 9871 6055 9877
rect 6822 9868 6828 9920
rect 6880 9908 6886 9920
rect 7208 9917 7236 9948
rect 7392 9948 7788 9976
rect 8113 9979 8171 9985
rect 7392 9917 7420 9948
rect 8113 9945 8125 9979
rect 8159 9976 8171 9979
rect 10054 9979 10112 9985
rect 10054 9976 10066 9979
rect 8159 9948 10066 9976
rect 8159 9945 8171 9948
rect 8113 9939 8171 9945
rect 10054 9945 10066 9948
rect 10100 9945 10112 9979
rect 10054 9939 10112 9945
rect 10796 9976 10824 10016
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11149 10047 11207 10053
rect 11149 10044 11161 10047
rect 11112 10016 11161 10044
rect 11112 10004 11118 10016
rect 11149 10013 11161 10016
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 11296 10016 11437 10044
rect 11296 10004 11302 10016
rect 11425 10013 11437 10016
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11606 10004 11612 10056
rect 11664 10004 11670 10056
rect 11790 10004 11796 10056
rect 11848 10004 11854 10056
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 12158 10044 12164 10056
rect 12023 10016 12164 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 12158 10004 12164 10016
rect 12216 10044 12222 10056
rect 12618 10044 12624 10056
rect 12216 10016 12624 10044
rect 12216 10004 12222 10016
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 12710 10004 12716 10056
rect 12768 10004 12774 10056
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10044 12863 10047
rect 12986 10044 12992 10056
rect 12851 10016 12992 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10013 13231 10047
rect 13173 10010 13231 10013
rect 13096 10007 13231 10010
rect 11333 9979 11391 9985
rect 11333 9976 11345 9979
rect 10796 9948 11345 9976
rect 7101 9911 7159 9917
rect 7101 9908 7113 9911
rect 6880 9880 7113 9908
rect 6880 9868 6886 9880
rect 7101 9877 7113 9880
rect 7147 9877 7159 9911
rect 7101 9871 7159 9877
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9877 7251 9911
rect 7193 9871 7251 9877
rect 7377 9911 7435 9917
rect 7377 9877 7389 9911
rect 7423 9877 7435 9911
rect 7377 9871 7435 9877
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10796 9908 10824 9948
rect 11333 9945 11345 9948
rect 11379 9945 11391 9979
rect 11333 9939 11391 9945
rect 13096 9982 13216 10007
rect 13446 10004 13452 10056
rect 13504 10004 13510 10056
rect 13817 10047 13875 10053
rect 13817 10013 13829 10047
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 9732 9880 10824 9908
rect 9732 9868 9738 9880
rect 12894 9868 12900 9920
rect 12952 9868 12958 9920
rect 13096 9917 13124 9982
rect 13832 9976 13860 10007
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 13964 10016 15025 10044
rect 13964 10004 13970 10016
rect 15013 10013 15025 10016
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 15102 10004 15108 10056
rect 15160 10004 15166 10056
rect 15194 10004 15200 10056
rect 15252 10004 15258 10056
rect 15304 10044 15332 10152
rect 15930 10072 15936 10124
rect 15988 10112 15994 10124
rect 16206 10112 16212 10124
rect 15988 10084 16212 10112
rect 15988 10072 15994 10084
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 16465 10047 16523 10053
rect 16465 10044 16477 10047
rect 15304 10016 16477 10044
rect 16465 10013 16477 10016
rect 16511 10013 16523 10047
rect 16465 10007 16523 10013
rect 15120 9976 15148 10004
rect 13832 9948 15148 9976
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9877 13139 9911
rect 13081 9871 13139 9877
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 13228 9880 13277 9908
rect 13228 9868 13234 9880
rect 13265 9877 13277 9880
rect 13311 9908 13323 9911
rect 13725 9911 13783 9917
rect 13725 9908 13737 9911
rect 13311 9880 13737 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 13725 9877 13737 9880
rect 13771 9877 13783 9911
rect 13725 9871 13783 9877
rect 15105 9911 15163 9917
rect 15105 9877 15117 9911
rect 15151 9908 15163 9911
rect 16022 9908 16028 9920
rect 15151 9880 16028 9908
rect 15151 9877 15163 9880
rect 15105 9871 15163 9877
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 1104 9818 18124 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 18124 9818
rect 1104 9744 18124 9766
rect 1762 9664 1768 9716
rect 1820 9704 1826 9716
rect 3237 9707 3295 9713
rect 3237 9704 3249 9707
rect 1820 9676 3249 9704
rect 1820 9664 1826 9676
rect 3237 9673 3249 9676
rect 3283 9673 3295 9707
rect 3237 9667 3295 9673
rect 3878 9664 3884 9716
rect 3936 9664 3942 9716
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 5721 9707 5779 9713
rect 5721 9704 5733 9707
rect 5684 9676 5733 9704
rect 5684 9664 5690 9676
rect 5721 9673 5733 9676
rect 5767 9673 5779 9707
rect 5721 9667 5779 9673
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 6730 9704 6736 9716
rect 5868 9676 6736 9704
rect 5868 9664 5874 9676
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 8389 9707 8447 9713
rect 8389 9673 8401 9707
rect 8435 9704 8447 9707
rect 8478 9704 8484 9716
rect 8435 9676 8484 9704
rect 8435 9673 8447 9676
rect 8389 9667 8447 9673
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 13081 9707 13139 9713
rect 13081 9704 13093 9707
rect 12768 9676 13093 9704
rect 12768 9664 12774 9676
rect 13081 9673 13093 9676
rect 13127 9673 13139 9707
rect 13081 9667 13139 9673
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 1857 9639 1915 9645
rect 1857 9636 1869 9639
rect 1728 9608 1869 9636
rect 1728 9596 1734 9608
rect 1857 9605 1869 9608
rect 1903 9605 1915 9639
rect 1857 9599 1915 9605
rect 2041 9639 2099 9645
rect 2041 9605 2053 9639
rect 2087 9636 2099 9639
rect 2501 9639 2559 9645
rect 2501 9636 2513 9639
rect 2087 9608 2513 9636
rect 2087 9605 2099 9608
rect 2041 9599 2099 9605
rect 2501 9605 2513 9608
rect 2547 9605 2559 9639
rect 6822 9636 6828 9648
rect 2501 9599 2559 9605
rect 5644 9608 6828 9636
rect 1765 9571 1823 9577
rect 1765 9568 1777 9571
rect 1504 9540 1777 9568
rect 1504 9364 1532 9540
rect 1765 9537 1777 9540
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 2130 9528 2136 9580
rect 2188 9577 2194 9580
rect 2188 9568 2197 9577
rect 2188 9540 2233 9568
rect 2188 9531 2197 9540
rect 2188 9528 2194 9531
rect 2958 9528 2964 9580
rect 3016 9568 3022 9580
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 3016 9540 3617 9568
rect 3016 9528 3022 9540
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 5534 9568 5540 9580
rect 4111 9540 5540 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 5644 9577 5672 9608
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 12161 9639 12219 9645
rect 12161 9605 12173 9639
rect 12207 9636 12219 9639
rect 12207 9608 13032 9636
rect 12207 9605 12219 9608
rect 12161 9599 12219 9605
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5960 9540 6009 9568
rect 5960 9528 5966 9540
rect 5997 9537 6009 9540
rect 6043 9537 6055 9571
rect 7190 9568 7196 9580
rect 5997 9531 6055 9537
rect 6104 9540 7196 9568
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 3418 9500 3424 9512
rect 3108 9472 3424 9500
rect 3108 9460 3114 9472
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 1578 9392 1584 9444
rect 1636 9432 1642 9444
rect 2041 9435 2099 9441
rect 2041 9432 2053 9435
rect 1636 9404 2053 9432
rect 1636 9392 1642 9404
rect 2041 9401 2053 9404
rect 2087 9401 2099 9435
rect 2041 9395 2099 9401
rect 2317 9435 2375 9441
rect 2317 9401 2329 9435
rect 2363 9432 2375 9435
rect 3528 9432 3556 9463
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 3752 9472 4169 9500
rect 3752 9460 3758 9472
rect 4157 9469 4169 9472
rect 4203 9469 4215 9503
rect 4157 9463 4215 9469
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9500 4307 9503
rect 4614 9500 4620 9512
rect 4295 9472 4620 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 6104 9432 6132 9540
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 8110 9528 8116 9580
rect 8168 9528 8174 9580
rect 8202 9528 8208 9580
rect 8260 9528 8266 9580
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 8352 9540 8401 9568
rect 8352 9528 8358 9540
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 9674 9528 9680 9580
rect 9732 9528 9738 9580
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 8478 9500 8484 9512
rect 6604 9472 8484 9500
rect 6604 9460 6610 9472
rect 8478 9460 8484 9472
rect 8536 9500 8542 9512
rect 9585 9503 9643 9509
rect 9585 9500 9597 9503
rect 8536 9472 9597 9500
rect 8536 9460 8542 9472
rect 9585 9469 9597 9472
rect 9631 9469 9643 9503
rect 9968 9500 9996 9531
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9568 10931 9571
rect 11054 9568 11060 9580
rect 10919 9540 11060 9568
rect 10919 9537 10931 9540
rect 10873 9531 10931 9537
rect 10888 9500 10916 9531
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 11146 9528 11152 9580
rect 11204 9528 11210 9580
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11606 9568 11612 9580
rect 11379 9540 11612 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 9968 9472 10916 9500
rect 9585 9463 9643 9469
rect 12158 9460 12164 9512
rect 12216 9460 12222 9512
rect 12452 9500 12480 9531
rect 12618 9528 12624 9580
rect 12676 9528 12682 9580
rect 12894 9528 12900 9580
rect 12952 9528 12958 9580
rect 12710 9500 12716 9512
rect 12452 9472 12716 9500
rect 12710 9460 12716 9472
rect 12768 9500 12774 9512
rect 13004 9500 13032 9608
rect 13096 9568 13124 9667
rect 13262 9664 13268 9716
rect 13320 9664 13326 9716
rect 13354 9664 13360 9716
rect 13412 9664 13418 9716
rect 14550 9664 14556 9716
rect 14608 9664 14614 9716
rect 14705 9639 14763 9645
rect 14705 9636 14717 9639
rect 14200 9608 14717 9636
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 13096 9540 13185 9568
rect 13173 9537 13185 9540
rect 13219 9537 13231 9571
rect 13906 9568 13912 9580
rect 13173 9531 13231 9537
rect 13372 9540 13912 9568
rect 13372 9500 13400 9540
rect 13906 9528 13912 9540
rect 13964 9528 13970 9580
rect 14200 9577 14228 9608
rect 14705 9605 14717 9608
rect 14751 9605 14763 9639
rect 14705 9599 14763 9605
rect 14918 9596 14924 9648
rect 14976 9636 14982 9648
rect 14976 9608 17540 9636
rect 14976 9596 14982 9608
rect 14185 9571 14243 9577
rect 14185 9537 14197 9571
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 14936 9568 14964 9596
rect 14507 9540 14964 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 12768 9472 12940 9500
rect 13004 9472 13400 9500
rect 12768 9460 12774 9472
rect 2363 9404 6132 9432
rect 6825 9435 6883 9441
rect 2363 9401 2375 9404
rect 2317 9395 2375 9401
rect 6825 9401 6837 9435
rect 6871 9432 6883 9435
rect 6914 9432 6920 9444
rect 6871 9404 6920 9432
rect 6871 9401 6883 9404
rect 6825 9395 6883 9401
rect 1946 9364 1952 9376
rect 1504 9336 1952 9364
rect 1946 9324 1952 9336
rect 2004 9364 2010 9376
rect 2332 9364 2360 9395
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 11057 9435 11115 9441
rect 11057 9401 11069 9435
rect 11103 9432 11115 9435
rect 11790 9432 11796 9444
rect 11103 9404 11796 9432
rect 11103 9401 11115 9404
rect 11057 9395 11115 9401
rect 11790 9392 11796 9404
rect 11848 9432 11854 9444
rect 12345 9435 12403 9441
rect 12345 9432 12357 9435
rect 11848 9404 12357 9432
rect 11848 9392 11854 9404
rect 12345 9401 12357 9404
rect 12391 9401 12403 9435
rect 12345 9395 12403 9401
rect 12805 9435 12863 9441
rect 12805 9401 12817 9435
rect 12851 9401 12863 9435
rect 12912 9432 12940 9472
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 14200 9500 14228 9531
rect 13596 9472 14228 9500
rect 14384 9500 14412 9531
rect 15102 9528 15108 9580
rect 15160 9528 15166 9580
rect 15764 9577 15792 9608
rect 17512 9580 17540 9608
rect 15749 9571 15807 9577
rect 15749 9537 15761 9571
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9537 16175 9571
rect 16117 9531 16175 9537
rect 16132 9500 16160 9531
rect 16206 9528 16212 9580
rect 16264 9528 16270 9580
rect 17494 9528 17500 9580
rect 17552 9528 17558 9580
rect 17402 9500 17408 9512
rect 14384 9472 14780 9500
rect 13596 9460 13602 9472
rect 14277 9435 14335 9441
rect 14277 9432 14289 9435
rect 12912 9404 14289 9432
rect 12805 9395 12863 9401
rect 14277 9401 14289 9404
rect 14323 9401 14335 9435
rect 14277 9395 14335 9401
rect 14752 9432 14780 9472
rect 16132 9472 17408 9500
rect 16132 9432 16160 9472
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 14752 9404 16160 9432
rect 2004 9336 2360 9364
rect 5905 9367 5963 9373
rect 2004 9324 2010 9336
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 6362 9364 6368 9376
rect 5951 9336 6368 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 12250 9364 12256 9376
rect 11664 9336 12256 9364
rect 11664 9324 11670 9336
rect 12250 9324 12256 9336
rect 12308 9364 12314 9376
rect 12820 9364 12848 9395
rect 12308 9336 12848 9364
rect 12308 9324 12314 9336
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 13044 9336 13277 9364
rect 13044 9324 13050 9336
rect 13265 9333 13277 9336
rect 13311 9333 13323 9367
rect 13265 9327 13323 9333
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 14752 9373 14780 9404
rect 17678 9392 17684 9444
rect 17736 9392 17742 9444
rect 14737 9367 14795 9373
rect 14737 9364 14749 9367
rect 14700 9336 14749 9364
rect 14700 9324 14706 9336
rect 14737 9333 14749 9336
rect 14783 9333 14795 9367
rect 14737 9327 14795 9333
rect 14826 9324 14832 9376
rect 14884 9364 14890 9376
rect 15010 9364 15016 9376
rect 14884 9336 15016 9364
rect 14884 9324 14890 9336
rect 15010 9324 15016 9336
rect 15068 9364 15074 9376
rect 15105 9367 15163 9373
rect 15105 9364 15117 9367
rect 15068 9336 15117 9364
rect 15068 9324 15074 9336
rect 15105 9333 15117 9336
rect 15151 9333 15163 9367
rect 15105 9327 15163 9333
rect 1104 9274 18124 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 18124 9274
rect 1104 9200 18124 9222
rect 1578 9120 1584 9172
rect 1636 9160 1642 9172
rect 2958 9160 2964 9172
rect 1636 9132 2964 9160
rect 1636 9120 1642 9132
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 6362 9120 6368 9172
rect 6420 9120 6426 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 10318 9160 10324 9172
rect 6880 9132 10324 9160
rect 6880 9120 6886 9132
rect 5902 9052 5908 9104
rect 5960 9092 5966 9104
rect 6454 9092 6460 9104
rect 5960 9064 6460 9092
rect 5960 9052 5966 9064
rect 6454 9052 6460 9064
rect 6512 9092 6518 9104
rect 7650 9092 7656 9104
rect 6512 9064 7656 9092
rect 6512 9052 6518 9064
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 5721 9027 5779 9033
rect 5721 8993 5733 9027
rect 5767 9024 5779 9027
rect 6546 9024 6552 9036
rect 5767 8996 6552 9024
rect 5767 8993 5779 8996
rect 5721 8987 5779 8993
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 8312 9033 8340 9132
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 12618 9120 12624 9172
rect 12676 9120 12682 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 12860 9132 12909 9160
rect 12860 9120 12866 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 15194 9120 15200 9172
rect 15252 9120 15258 9172
rect 17313 9163 17371 9169
rect 17313 9129 17325 9163
rect 17359 9160 17371 9163
rect 17494 9160 17500 9172
rect 17359 9132 17500 9160
rect 17359 9129 17371 9132
rect 17313 9123 17371 9129
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 9493 9095 9551 9101
rect 9493 9061 9505 9095
rect 9539 9061 9551 9095
rect 12636 9092 12664 9120
rect 14458 9092 14464 9104
rect 12636 9064 14464 9092
rect 9493 9055 9551 9061
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 8993 8355 9027
rect 8297 8987 8355 8993
rect 8478 8984 8484 9036
rect 8536 8984 8542 9036
rect 9508 9024 9536 9055
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 10502 9024 10508 9036
rect 9508 8996 10508 9024
rect 10502 8984 10508 8996
rect 10560 9024 10566 9036
rect 10560 8996 10732 9024
rect 10560 8984 10566 8996
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 6822 8956 6828 8968
rect 5951 8928 6828 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 9214 8956 9220 8968
rect 8619 8928 9220 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 6454 8897 6460 8900
rect 6181 8891 6239 8897
rect 6181 8857 6193 8891
rect 6227 8857 6239 8891
rect 6181 8851 6239 8857
rect 6397 8891 6460 8897
rect 6397 8857 6409 8891
rect 6443 8857 6460 8891
rect 6397 8851 6460 8857
rect 6089 8823 6147 8829
rect 6089 8789 6101 8823
rect 6135 8820 6147 8823
rect 6196 8820 6224 8851
rect 6454 8848 6460 8851
rect 6512 8848 6518 8900
rect 6730 8848 6736 8900
rect 6788 8888 6794 8900
rect 8404 8888 8432 8919
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9490 8916 9496 8968
rect 9548 8916 9554 8968
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 6788 8860 8432 8888
rect 6788 8848 6794 8860
rect 6135 8792 6224 8820
rect 6135 8789 6147 8792
rect 6089 8783 6147 8789
rect 6546 8780 6552 8832
rect 6604 8780 6610 8832
rect 7190 8780 7196 8832
rect 7248 8820 7254 8832
rect 8113 8823 8171 8829
rect 8113 8820 8125 8823
rect 7248 8792 8125 8820
rect 7248 8780 7254 8792
rect 8113 8789 8125 8792
rect 8159 8789 8171 8823
rect 8404 8820 8432 8860
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 9600 8888 9628 8919
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 10704 8965 10732 8996
rect 11422 8984 11428 9036
rect 11480 9024 11486 9036
rect 12621 9027 12679 9033
rect 12621 9024 12633 9027
rect 11480 8996 12633 9024
rect 11480 8984 11486 8996
rect 12621 8993 12633 8996
rect 12667 8993 12679 9027
rect 12621 8987 12679 8993
rect 12710 8984 12716 9036
rect 12768 8984 12774 9036
rect 15930 8984 15936 9036
rect 15988 8984 15994 9036
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 10284 8928 10425 8956
rect 10284 8916 10290 8928
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 12250 8916 12256 8968
rect 12308 8956 12314 8968
rect 12419 8959 12477 8965
rect 12419 8956 12431 8959
rect 12308 8928 12431 8956
rect 12308 8916 12314 8928
rect 12406 8925 12431 8928
rect 12465 8925 12477 8959
rect 12406 8919 12477 8925
rect 12535 8959 12593 8965
rect 12535 8925 12547 8959
rect 12581 8956 12593 8959
rect 12894 8956 12900 8968
rect 12581 8928 12900 8956
rect 12581 8925 12593 8928
rect 12535 8919 12593 8925
rect 9364 8860 9628 8888
rect 9364 8848 9370 8860
rect 9766 8848 9772 8900
rect 9824 8848 9830 8900
rect 10597 8891 10655 8897
rect 10597 8857 10609 8891
rect 10643 8888 10655 8891
rect 12406 8888 12434 8919
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 14550 8916 14556 8968
rect 14608 8916 14614 8968
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8956 14795 8959
rect 14826 8956 14832 8968
rect 14783 8928 14832 8956
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15013 8959 15071 8965
rect 15013 8956 15025 8959
rect 14976 8928 15025 8956
rect 14976 8916 14982 8928
rect 15013 8925 15025 8928
rect 15059 8925 15071 8959
rect 15013 8919 15071 8925
rect 16022 8916 16028 8968
rect 16080 8956 16086 8968
rect 16189 8959 16247 8965
rect 16189 8956 16201 8959
rect 16080 8928 16201 8956
rect 16080 8916 16086 8928
rect 16189 8925 16201 8928
rect 16235 8925 16247 8959
rect 16189 8919 16247 8925
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 14366 8888 14372 8900
rect 10643 8860 11468 8888
rect 12406 8860 14372 8888
rect 10643 8857 10655 8860
rect 10597 8851 10655 8857
rect 10873 8823 10931 8829
rect 10873 8820 10885 8823
rect 8404 8792 10885 8820
rect 8113 8783 8171 8789
rect 10873 8789 10885 8792
rect 10919 8789 10931 8823
rect 11440 8820 11468 8860
rect 14366 8848 14372 8860
rect 14424 8848 14430 8900
rect 17512 8888 17540 8919
rect 16224 8860 17540 8888
rect 16224 8832 16252 8860
rect 13354 8820 13360 8832
rect 11440 8792 13360 8820
rect 10873 8783 10931 8789
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 16206 8780 16212 8832
rect 16264 8780 16270 8832
rect 17678 8780 17684 8832
rect 17736 8780 17742 8832
rect 1104 8730 18124 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 18124 8730
rect 1104 8656 18124 8678
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7558 8616 7564 8628
rect 7515 8588 7564 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7558 8576 7564 8588
rect 7616 8616 7622 8628
rect 7616 8588 8156 8616
rect 7616 8576 7622 8588
rect 7653 8551 7711 8557
rect 7653 8517 7665 8551
rect 7699 8548 7711 8551
rect 8018 8548 8024 8560
rect 7699 8520 8024 8548
rect 7699 8517 7711 8520
rect 7653 8511 7711 8517
rect 8018 8508 8024 8520
rect 8076 8508 8082 8560
rect 8128 8548 8156 8588
rect 9766 8576 9772 8628
rect 9824 8616 9830 8628
rect 11149 8619 11207 8625
rect 11149 8616 11161 8619
rect 9824 8588 11161 8616
rect 9824 8576 9830 8588
rect 11149 8585 11161 8588
rect 11195 8616 11207 8619
rect 11422 8616 11428 8628
rect 11195 8588 11428 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 11532 8588 14136 8616
rect 10594 8548 10600 8560
rect 8128 8520 10600 8548
rect 10594 8508 10600 8520
rect 10652 8508 10658 8560
rect 11330 8548 11336 8560
rect 11072 8520 11336 8548
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 1946 8480 1952 8492
rect 1903 8452 1952 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8480 2283 8483
rect 3142 8480 3148 8492
rect 2271 8452 3148 8480
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 7374 8440 7380 8492
rect 7432 8440 7438 8492
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8480 7803 8483
rect 7926 8480 7932 8492
rect 7791 8452 7932 8480
rect 7791 8449 7803 8452
rect 7745 8443 7803 8449
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 11072 8489 11100 8520
rect 11330 8508 11336 8520
rect 11388 8548 11394 8560
rect 11532 8548 11560 8588
rect 11388 8520 11560 8548
rect 11793 8551 11851 8557
rect 11388 8508 11394 8520
rect 11793 8517 11805 8551
rect 11839 8548 11851 8551
rect 12250 8548 12256 8560
rect 11839 8520 12256 8548
rect 11839 8517 11851 8520
rect 11793 8511 11851 8517
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 14108 8489 14136 8588
rect 14366 8508 14372 8560
rect 14424 8548 14430 8560
rect 14424 8520 15056 8548
rect 14424 8508 14430 8520
rect 11609 8483 11667 8489
rect 11609 8480 11621 8483
rect 11204 8452 11621 8480
rect 11204 8440 11210 8452
rect 11609 8449 11621 8452
rect 11655 8480 11667 8483
rect 14093 8483 14151 8489
rect 11655 8452 12572 8480
rect 11655 8449 11667 8452
rect 11609 8443 11667 8449
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 5868 8384 8033 8412
rect 5868 8372 5874 8384
rect 8021 8381 8033 8384
rect 8067 8412 8079 8415
rect 9214 8412 9220 8424
rect 8067 8384 9220 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 2038 8304 2044 8356
rect 2096 8304 2102 8356
rect 7653 8347 7711 8353
rect 7653 8313 7665 8347
rect 7699 8344 7711 8347
rect 7837 8347 7895 8353
rect 7837 8344 7849 8347
rect 7699 8316 7849 8344
rect 7699 8313 7711 8316
rect 7653 8307 7711 8313
rect 7837 8313 7849 8316
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 10321 8347 10379 8353
rect 10321 8344 10333 8347
rect 8168 8316 10333 8344
rect 8168 8304 8174 8316
rect 10321 8313 10333 8316
rect 10367 8344 10379 8347
rect 12250 8344 12256 8356
rect 10367 8316 12256 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 12250 8304 12256 8316
rect 12308 8304 12314 8356
rect 12544 8344 12572 8452
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14277 8483 14335 8489
rect 14277 8449 14289 8483
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 13538 8412 13544 8424
rect 12676 8384 13544 8412
rect 12676 8372 12682 8384
rect 13538 8372 13544 8384
rect 13596 8412 13602 8424
rect 14292 8412 14320 8443
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 14734 8440 14740 8492
rect 14792 8440 14798 8492
rect 15028 8489 15056 8520
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 17402 8440 17408 8492
rect 17460 8480 17466 8492
rect 17497 8483 17555 8489
rect 17497 8480 17509 8483
rect 17460 8452 17509 8480
rect 17460 8440 17466 8452
rect 17497 8449 17509 8452
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 15470 8412 15476 8424
rect 13596 8384 15476 8412
rect 13596 8372 13602 8384
rect 15470 8372 15476 8384
rect 15528 8412 15534 8424
rect 16206 8412 16212 8424
rect 15528 8384 16212 8412
rect 15528 8372 15534 8384
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 14734 8344 14740 8356
rect 12544 8316 14740 8344
rect 14734 8304 14740 8316
rect 14792 8304 14798 8356
rect 14826 8304 14832 8356
rect 14884 8304 14890 8356
rect 17678 8304 17684 8356
rect 17736 8304 17742 8356
rect 1486 8236 1492 8288
rect 1544 8276 1550 8288
rect 1673 8279 1731 8285
rect 1673 8276 1685 8279
rect 1544 8248 1685 8276
rect 1544 8236 1550 8248
rect 1673 8245 1685 8248
rect 1719 8276 1731 8279
rect 3326 8276 3332 8288
rect 1719 8248 3332 8276
rect 1719 8245 1731 8248
rect 1673 8239 1731 8245
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 7742 8236 7748 8288
rect 7800 8236 7806 8288
rect 11974 8236 11980 8288
rect 12032 8236 12038 8288
rect 1104 8186 18124 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 18124 8186
rect 1104 8112 18124 8134
rect 3142 8032 3148 8084
rect 3200 8032 3206 8084
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 5626 8072 5632 8084
rect 5491 8044 5632 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 7432 8044 9045 8072
rect 7432 8032 7438 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 9490 8032 9496 8084
rect 9548 8072 9554 8084
rect 11241 8075 11299 8081
rect 11241 8072 11253 8075
rect 9548 8044 11253 8072
rect 9548 8032 9554 8044
rect 11241 8041 11253 8044
rect 11287 8041 11299 8075
rect 11241 8035 11299 8041
rect 12618 8032 12624 8084
rect 12676 8032 12682 8084
rect 12986 8032 12992 8084
rect 13044 8032 13050 8084
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 3160 7936 3188 8032
rect 9398 8004 9404 8016
rect 9232 7976 9404 8004
rect 3605 7939 3663 7945
rect 3605 7936 3617 7939
rect 3160 7908 3617 7936
rect 3605 7905 3617 7908
rect 3651 7936 3663 7939
rect 6825 7939 6883 7945
rect 3651 7908 4200 7936
rect 3651 7905 3663 7908
rect 3605 7899 3663 7905
rect 1670 7828 1676 7880
rect 1728 7828 1734 7880
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7868 1823 7871
rect 1854 7868 1860 7880
rect 1811 7840 1860 7868
rect 1811 7837 1823 7840
rect 1765 7831 1823 7837
rect 1854 7828 1860 7840
rect 1912 7828 1918 7880
rect 3418 7868 3424 7880
rect 1964 7840 3424 7868
rect 1394 7760 1400 7812
rect 1452 7800 1458 7812
rect 1964 7800 1992 7840
rect 3418 7828 3424 7840
rect 3476 7868 3482 7880
rect 4172 7877 4200 7908
rect 6825 7905 6837 7939
rect 6871 7936 6883 7939
rect 6914 7936 6920 7948
rect 6871 7908 6920 7936
rect 6871 7905 6883 7908
rect 6825 7899 6883 7905
rect 6914 7896 6920 7908
rect 6972 7936 6978 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 6972 7908 7205 7936
rect 6972 7896 6978 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3476 7840 3801 7868
rect 3476 7828 3482 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4706 7828 4712 7880
rect 4764 7828 4770 7880
rect 4798 7828 4804 7880
rect 4856 7868 4862 7880
rect 5077 7871 5135 7877
rect 5077 7868 5089 7871
rect 4856 7840 5089 7868
rect 4856 7828 4862 7840
rect 5077 7837 5089 7840
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 6546 7828 6552 7880
rect 6604 7877 6610 7880
rect 6604 7868 6616 7877
rect 7460 7871 7518 7877
rect 6604 7840 6649 7868
rect 6604 7831 6616 7840
rect 7460 7837 7472 7871
rect 7506 7868 7518 7871
rect 7742 7868 7748 7880
rect 7506 7840 7748 7868
rect 7506 7837 7518 7840
rect 7460 7831 7518 7837
rect 6604 7828 6610 7831
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 9232 7877 9260 7976
rect 9398 7964 9404 7976
rect 9456 8004 9462 8016
rect 11057 8007 11115 8013
rect 11057 8004 11069 8007
rect 9456 7976 11069 8004
rect 9456 7964 9462 7976
rect 11057 7973 11069 7976
rect 11103 7973 11115 8007
rect 11057 7967 11115 7973
rect 12526 7964 12532 8016
rect 12584 8004 12590 8016
rect 14737 8007 14795 8013
rect 12584 7976 14596 8004
rect 12584 7964 12590 7976
rect 10137 7939 10195 7945
rect 9324 7908 10088 7936
rect 9324 7880 9352 7908
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9548 7840 9597 7868
rect 9548 7828 9554 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 1452 7772 1992 7800
rect 2032 7803 2090 7809
rect 1452 7760 1458 7772
rect 2032 7769 2044 7803
rect 2078 7800 2090 7803
rect 2314 7800 2320 7812
rect 2078 7772 2320 7800
rect 2078 7769 2090 7772
rect 2032 7763 2090 7769
rect 2314 7760 2320 7772
rect 2372 7760 2378 7812
rect 4985 7803 5043 7809
rect 4985 7769 4997 7803
rect 5031 7800 5043 7803
rect 9324 7800 9352 7828
rect 5031 7772 9352 7800
rect 9600 7800 9628 7831
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 10060 7868 10088 7908
rect 10137 7905 10149 7939
rect 10183 7936 10195 7939
rect 10226 7936 10232 7948
rect 10183 7908 10232 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 10336 7908 11345 7936
rect 10060 7864 10272 7868
rect 10336 7864 10364 7908
rect 10704 7877 10732 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 11422 7896 11428 7948
rect 11480 7896 11486 7948
rect 12066 7896 12072 7948
rect 12124 7936 12130 7948
rect 12124 7908 12388 7936
rect 12124 7896 12130 7908
rect 10060 7840 10364 7864
rect 10244 7836 10364 7840
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 11440 7868 11468 7896
rect 12360 7877 12388 7908
rect 12986 7896 12992 7948
rect 13044 7936 13050 7948
rect 14568 7936 14596 7976
rect 14737 7973 14749 8007
rect 14783 8004 14795 8007
rect 16577 8007 16635 8013
rect 14783 7976 15240 8004
rect 14783 7973 14795 7976
rect 14737 7967 14795 7973
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 13044 7908 14504 7936
rect 14568 7908 14841 7936
rect 13044 7896 13050 7908
rect 14476 7877 14504 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 15212 7936 15240 7976
rect 16577 7973 16589 8007
rect 16623 7973 16635 8007
rect 16577 7967 16635 7973
rect 16592 7936 16620 7967
rect 17402 7936 17408 7948
rect 15212 7908 15332 7936
rect 16592 7908 17408 7936
rect 14829 7899 14887 7905
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11440 7840 12173 7868
rect 10689 7831 10747 7837
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7868 12403 7871
rect 14461 7871 14519 7877
rect 12391 7840 14412 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 10428 7800 10456 7831
rect 9600 7772 10456 7800
rect 5031 7769 5043 7772
rect 4985 7763 5043 7769
rect 10962 7760 10968 7812
rect 11020 7800 11026 7812
rect 11057 7803 11115 7809
rect 11057 7800 11069 7803
rect 11020 7772 11069 7800
rect 11020 7760 11026 7772
rect 11057 7769 11069 7772
rect 11103 7769 11115 7803
rect 12805 7803 12863 7809
rect 12805 7800 12817 7803
rect 11057 7763 11115 7769
rect 12452 7772 12817 7800
rect 842 7692 848 7744
rect 900 7732 906 7744
rect 1489 7735 1547 7741
rect 1489 7732 1501 7735
rect 900 7704 1501 7732
rect 900 7692 906 7704
rect 1489 7701 1501 7704
rect 1535 7701 1547 7735
rect 1489 7695 1547 7701
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 3510 7732 3516 7744
rect 3283 7704 3516 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 8573 7735 8631 7741
rect 8573 7732 8585 7735
rect 8076 7704 8585 7732
rect 8076 7692 8082 7704
rect 8573 7701 8585 7704
rect 8619 7701 8631 7735
rect 8573 7695 8631 7701
rect 10410 7692 10416 7744
rect 10468 7732 10474 7744
rect 12452 7741 12480 7772
rect 12805 7769 12817 7772
rect 12851 7769 12863 7803
rect 14384 7800 14412 7840
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14550 7828 14556 7880
rect 14608 7868 14614 7880
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14608 7840 15117 7868
rect 14608 7828 14614 7840
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15194 7828 15200 7880
rect 15252 7828 15258 7880
rect 15304 7868 15332 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 15453 7871 15511 7877
rect 15453 7868 15465 7871
rect 15304 7840 15465 7868
rect 15453 7837 15465 7840
rect 15499 7837 15511 7871
rect 15453 7831 15511 7837
rect 14568 7800 14596 7828
rect 14384 7772 14596 7800
rect 14737 7803 14795 7809
rect 12805 7763 12863 7769
rect 14737 7769 14749 7803
rect 14783 7800 14795 7803
rect 14829 7803 14887 7809
rect 14829 7800 14841 7803
rect 14783 7772 14841 7800
rect 14783 7769 14795 7772
rect 14737 7763 14795 7769
rect 14829 7769 14841 7772
rect 14875 7769 14887 7803
rect 14829 7763 14887 7769
rect 10689 7735 10747 7741
rect 10689 7732 10701 7735
rect 10468 7704 10701 7732
rect 10468 7692 10474 7704
rect 10689 7701 10701 7704
rect 10735 7701 10747 7735
rect 10689 7695 10747 7701
rect 12437 7735 12495 7741
rect 12437 7701 12449 7735
rect 12483 7701 12495 7735
rect 12437 7695 12495 7701
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 13005 7735 13063 7741
rect 13005 7732 13017 7735
rect 12584 7704 13017 7732
rect 12584 7692 12590 7704
rect 13005 7701 13017 7704
rect 13051 7701 13063 7735
rect 13005 7695 13063 7701
rect 13173 7735 13231 7741
rect 13173 7701 13185 7735
rect 13219 7732 13231 7735
rect 14182 7732 14188 7744
rect 13219 7704 14188 7732
rect 13219 7701 13231 7704
rect 13173 7695 13231 7701
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 14553 7735 14611 7741
rect 14553 7701 14565 7735
rect 14599 7732 14611 7735
rect 15746 7732 15752 7744
rect 14599 7704 15752 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 16758 7692 16764 7744
rect 16816 7692 16822 7744
rect 1104 7642 18124 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 18124 7642
rect 1104 7568 18124 7590
rect 1486 7488 1492 7540
rect 1544 7488 1550 7540
rect 2314 7488 2320 7540
rect 2372 7488 2378 7540
rect 4706 7488 4712 7540
rect 4764 7528 4770 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 4764 7500 5549 7528
rect 4764 7488 4770 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 5537 7491 5595 7497
rect 5810 7488 5816 7540
rect 5868 7488 5874 7540
rect 7926 7488 7932 7540
rect 7984 7488 7990 7540
rect 15470 7488 15476 7540
rect 15528 7488 15534 7540
rect 15746 7488 15752 7540
rect 15804 7488 15810 7540
rect 1854 7420 1860 7472
rect 1912 7460 1918 7472
rect 6914 7460 6920 7472
rect 1912 7432 6920 7460
rect 1912 7420 1918 7432
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 1765 7395 1823 7401
rect 1765 7392 1777 7395
rect 1688 7364 1777 7392
rect 1578 7284 1584 7336
rect 1636 7284 1642 7336
rect 1688 7188 1716 7364
rect 1765 7361 1777 7364
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 2130 7352 2136 7404
rect 2188 7352 2194 7404
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2455 7364 3280 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2240 7324 2268 7355
rect 1780 7296 2268 7324
rect 1780 7265 1808 7296
rect 3142 7284 3148 7336
rect 3200 7284 3206 7336
rect 3252 7333 3280 7364
rect 3326 7352 3332 7404
rect 3384 7392 3390 7404
rect 3421 7395 3479 7401
rect 3421 7392 3433 7395
rect 3384 7364 3433 7392
rect 3384 7352 3390 7364
rect 3421 7361 3433 7364
rect 3467 7361 3479 7395
rect 3421 7355 3479 7361
rect 3510 7352 3516 7404
rect 3568 7352 3574 7404
rect 3602 7352 3608 7404
rect 3660 7352 3666 7404
rect 4172 7401 4200 7432
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 7558 7420 7564 7472
rect 7616 7420 7622 7472
rect 7777 7463 7835 7469
rect 7777 7429 7789 7463
rect 7823 7460 7835 7463
rect 10137 7463 10195 7469
rect 7823 7432 7972 7460
rect 7823 7429 7835 7432
rect 7777 7423 7835 7429
rect 7944 7404 7972 7432
rect 10137 7429 10149 7463
rect 10183 7460 10195 7463
rect 10686 7460 10692 7472
rect 10183 7432 10692 7460
rect 10183 7429 10195 7432
rect 10137 7423 10195 7429
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 12066 7460 12072 7472
rect 11808 7432 12072 7460
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4424 7395 4482 7401
rect 4424 7361 4436 7395
rect 4470 7392 4482 7395
rect 4706 7392 4712 7404
rect 4470 7364 4712 7392
rect 4470 7361 4482 7364
rect 4424 7355 4482 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 5902 7392 5908 7404
rect 5767 7364 5908 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 7926 7352 7932 7404
rect 7984 7352 7990 7404
rect 9858 7352 9864 7404
rect 9916 7352 9922 7404
rect 9950 7352 9956 7404
rect 10008 7352 10014 7404
rect 10318 7352 10324 7404
rect 10376 7352 10382 7404
rect 10410 7352 10416 7404
rect 10468 7392 10474 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 10468 7364 10517 7392
rect 10468 7352 10474 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7392 10655 7395
rect 11330 7392 11336 7404
rect 10643 7364 11336 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 11808 7401 11836 7432
rect 12066 7420 12072 7432
rect 12124 7420 12130 7472
rect 12250 7420 12256 7472
rect 12308 7420 12314 7472
rect 15194 7460 15200 7472
rect 14108 7432 15200 7460
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 11974 7352 11980 7404
rect 12032 7352 12038 7404
rect 12802 7352 12808 7404
rect 12860 7392 12866 7404
rect 14108 7401 14136 7432
rect 15194 7420 15200 7432
rect 15252 7420 15258 7472
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 12860 7364 14013 7392
rect 12860 7352 12866 7364
rect 14001 7361 14013 7364
rect 14047 7392 14059 7395
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 14047 7364 14105 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 14349 7395 14407 7401
rect 14349 7392 14361 7395
rect 14240 7364 14361 7392
rect 14240 7352 14246 7364
rect 14349 7361 14361 7364
rect 14395 7361 14407 7395
rect 14349 7355 14407 7361
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7392 15899 7395
rect 16758 7392 16764 7404
rect 15887 7364 16764 7392
rect 15887 7361 15899 7364
rect 15841 7355 15899 7361
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7293 3295 7327
rect 3237 7287 3295 7293
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 9876 7324 9904 7352
rect 10226 7324 10232 7336
rect 3752 7296 4200 7324
rect 9876 7296 10232 7324
rect 3752 7284 3758 7296
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7225 1823 7259
rect 2501 7259 2559 7265
rect 2501 7256 2513 7259
rect 1765 7219 1823 7225
rect 1872 7228 2513 7256
rect 1872 7188 1900 7228
rect 2501 7225 2513 7228
rect 2547 7225 2559 7259
rect 2501 7219 2559 7225
rect 1688 7160 1900 7188
rect 1946 7148 1952 7200
rect 2004 7148 2010 7200
rect 4172 7188 4200 7296
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 5810 7188 5816 7200
rect 4172 7160 5816 7188
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 7558 7188 7564 7200
rect 7432 7160 7564 7188
rect 7432 7148 7438 7160
rect 7558 7148 7564 7160
rect 7616 7188 7622 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 7616 7160 7757 7188
rect 7616 7148 7622 7160
rect 7745 7157 7757 7160
rect 7791 7157 7803 7191
rect 7745 7151 7803 7157
rect 10597 7191 10655 7197
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 10643 7160 11529 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 11606 7148 11612 7200
rect 11664 7188 11670 7200
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11664 7160 11805 7188
rect 11664 7148 11670 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 11793 7151 11851 7157
rect 1104 7098 18124 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 18124 7098
rect 1104 7024 18124 7046
rect 4525 6987 4583 6993
rect 4525 6953 4537 6987
rect 4571 6984 4583 6987
rect 4706 6984 4712 6996
rect 4571 6956 4712 6984
rect 4571 6953 4583 6956
rect 4525 6947 4583 6953
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 10137 6987 10195 6993
rect 10137 6953 10149 6987
rect 10183 6984 10195 6987
rect 10318 6984 10324 6996
rect 10183 6956 10324 6984
rect 10183 6953 10195 6956
rect 10137 6947 10195 6953
rect 10318 6944 10324 6956
rect 10376 6944 10382 6996
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 4614 6916 4620 6928
rect 4212 6888 4620 6916
rect 4212 6876 4218 6888
rect 4614 6876 4620 6888
rect 4672 6876 4678 6928
rect 5902 6916 5908 6928
rect 5460 6888 5908 6916
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 2774 6848 2780 6860
rect 1636 6820 2780 6848
rect 1636 6808 1642 6820
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 3602 6808 3608 6860
rect 3660 6848 3666 6860
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3660 6820 3985 6848
rect 3660 6808 3666 6820
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 4120 6820 4660 6848
rect 4120 6808 4126 6820
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 2130 6780 2136 6792
rect 1903 6752 2136 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 2455 6752 2513 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2501 6749 2513 6752
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 3326 6780 3332 6792
rect 3016 6752 3332 6780
rect 3016 6740 3022 6752
rect 3326 6740 3332 6752
rect 3384 6780 3390 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3384 6752 3801 6780
rect 3384 6740 3390 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 4154 6740 4160 6792
rect 4212 6740 4218 6792
rect 4632 6789 4660 6820
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6780 4859 6783
rect 5460 6780 5488 6888
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 11793 6919 11851 6925
rect 11793 6885 11805 6919
rect 11839 6916 11851 6919
rect 12069 6919 12127 6925
rect 12069 6916 12081 6919
rect 11839 6888 12081 6916
rect 11839 6885 11851 6888
rect 11793 6879 11851 6885
rect 12069 6885 12081 6888
rect 12115 6885 12127 6919
rect 12069 6879 12127 6885
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 10962 6848 10968 6860
rect 9723 6820 10180 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 4847 6752 5488 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 4356 6712 4384 6743
rect 4080 6684 4384 6712
rect 4540 6712 4568 6743
rect 9582 6740 9588 6792
rect 9640 6740 9646 6792
rect 10152 6789 10180 6820
rect 10336 6820 10968 6848
rect 10336 6792 10364 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11330 6808 11336 6860
rect 11388 6848 11394 6860
rect 11388 6820 11744 6848
rect 11388 6808 11394 6820
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 4709 6715 4767 6721
rect 4709 6712 4721 6715
rect 4540 6684 4721 6712
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2593 6647 2651 6653
rect 2593 6644 2605 6647
rect 2004 6616 2605 6644
rect 2004 6604 2010 6616
rect 2593 6613 2605 6616
rect 2639 6613 2651 6647
rect 2593 6607 2651 6613
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 4080 6653 4108 6684
rect 4709 6681 4721 6684
rect 4755 6681 4767 6715
rect 4709 6675 4767 6681
rect 6641 6715 6699 6721
rect 6641 6681 6653 6715
rect 6687 6712 6699 6715
rect 6914 6712 6920 6724
rect 6687 6684 6920 6712
rect 6687 6681 6699 6684
rect 6641 6675 6699 6681
rect 6914 6672 6920 6684
rect 6972 6672 6978 6724
rect 8570 6672 8576 6724
rect 8628 6712 8634 6724
rect 9784 6712 9812 6743
rect 10318 6740 10324 6792
rect 10376 6740 10382 6792
rect 10410 6740 10416 6792
rect 10468 6780 10474 6792
rect 10468 6752 10548 6780
rect 10468 6740 10474 6752
rect 10520 6712 10548 6752
rect 10594 6740 10600 6792
rect 10652 6740 10658 6792
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 11606 6780 11612 6792
rect 10827 6752 11612 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 11716 6789 11744 6820
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 12032 6820 12572 6848
rect 12032 6808 12038 6820
rect 11701 6783 11759 6789
rect 11701 6749 11713 6783
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 11793 6783 11851 6789
rect 11793 6749 11805 6783
rect 11839 6780 11851 6783
rect 11882 6780 11888 6792
rect 11839 6752 11888 6780
rect 11839 6749 11851 6752
rect 11793 6743 11851 6749
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 12066 6740 12072 6792
rect 12124 6780 12130 6792
rect 12544 6789 12572 6820
rect 12345 6783 12403 6789
rect 12345 6780 12357 6783
rect 12124 6752 12357 6780
rect 12124 6740 12130 6752
rect 12345 6749 12357 6752
rect 12391 6749 12403 6783
rect 12345 6743 12403 6749
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12802 6740 12808 6792
rect 12860 6740 12866 6792
rect 11517 6715 11575 6721
rect 11517 6712 11529 6715
rect 8628 6684 10456 6712
rect 10520 6684 11529 6712
rect 8628 6672 8634 6684
rect 10428 6656 10456 6684
rect 11517 6681 11529 6684
rect 11563 6681 11575 6715
rect 11517 6675 11575 6681
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3568 6616 3893 6644
rect 3568 6604 3574 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 3881 6607 3939 6613
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 10410 6604 10416 6656
rect 10468 6604 10474 6656
rect 10781 6647 10839 6653
rect 10781 6613 10793 6647
rect 10827 6644 10839 6647
rect 10870 6644 10876 6656
rect 10827 6616 10876 6644
rect 10827 6613 10839 6616
rect 10781 6607 10839 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 11532 6644 11560 6675
rect 12434 6672 12440 6724
rect 12492 6712 12498 6724
rect 12820 6712 12848 6740
rect 12492 6684 12848 6712
rect 12492 6672 12498 6684
rect 11606 6644 11612 6656
rect 11532 6616 11612 6644
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 12250 6604 12256 6656
rect 12308 6604 12314 6656
rect 1104 6554 18124 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 18124 6554
rect 1104 6480 18124 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 2130 6440 2136 6452
rect 1627 6412 2136 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 2130 6400 2136 6412
rect 2188 6440 2194 6452
rect 3221 6443 3279 6449
rect 2188 6412 2774 6440
rect 2188 6400 2194 6412
rect 2746 6372 2774 6412
rect 3221 6409 3233 6443
rect 3267 6440 3279 6443
rect 3510 6440 3516 6452
rect 3267 6412 3516 6440
rect 3267 6409 3279 6412
rect 3221 6403 3279 6409
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 9398 6400 9404 6452
rect 9456 6400 9462 6452
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 12526 6440 12532 6452
rect 10652 6412 12532 6440
rect 10652 6400 10658 6412
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 3421 6375 3479 6381
rect 3421 6372 3433 6375
rect 2746 6344 3433 6372
rect 3421 6341 3433 6344
rect 3467 6372 3479 6375
rect 4798 6372 4804 6384
rect 3467 6344 4804 6372
rect 3467 6341 3479 6344
rect 3421 6335 3479 6341
rect 4798 6332 4804 6344
rect 4856 6332 4862 6384
rect 8110 6332 8116 6384
rect 8168 6332 8174 6384
rect 9950 6372 9956 6384
rect 9048 6344 9956 6372
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2694 6307 2752 6313
rect 2694 6304 2706 6307
rect 2188 6276 2706 6304
rect 2188 6264 2194 6276
rect 2694 6273 2706 6276
rect 2740 6273 2752 6307
rect 2694 6267 2752 6273
rect 7926 6264 7932 6316
rect 7984 6304 7990 6316
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 7984 6276 8309 6304
rect 7984 6264 7990 6276
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 4614 6236 4620 6248
rect 3007 6208 4620 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 4614 6196 4620 6208
rect 4672 6196 4678 6248
rect 2976 6140 3280 6168
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 2976 6100 3004 6140
rect 1728 6072 3004 6100
rect 1728 6060 1734 6072
rect 3050 6060 3056 6112
rect 3108 6060 3114 6112
rect 3252 6109 3280 6140
rect 3602 6128 3608 6180
rect 3660 6168 3666 6180
rect 8312 6168 8340 6267
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 9048 6313 9076 6344
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 8772 6236 8800 6267
rect 9122 6264 9128 6316
rect 9180 6264 9186 6316
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9582 6304 9588 6316
rect 9355 6276 9588 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 8444 6208 8800 6236
rect 8444 6196 8450 6208
rect 9324 6168 9352 6267
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6304 9735 6307
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9723 6276 9781 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 10502 6264 10508 6316
rect 10560 6264 10566 6316
rect 10870 6264 10876 6316
rect 10928 6264 10934 6316
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6273 11115 6307
rect 11057 6267 11115 6273
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 9493 6199 9551 6205
rect 3660 6140 8248 6168
rect 8312 6140 9352 6168
rect 3660 6128 3666 6140
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6100 3295 6103
rect 3970 6100 3976 6112
rect 3283 6072 3976 6100
rect 3283 6069 3295 6072
rect 3237 6063 3295 6069
rect 3970 6060 3976 6072
rect 4028 6100 4034 6112
rect 4154 6100 4160 6112
rect 4028 6072 4160 6100
rect 4028 6060 4034 6072
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 6825 6103 6883 6109
rect 6825 6069 6837 6103
rect 6871 6100 6883 6103
rect 6914 6100 6920 6112
rect 6871 6072 6920 6100
rect 6871 6069 6883 6072
rect 6825 6063 6883 6069
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 8220 6100 8248 6140
rect 9030 6100 9036 6112
rect 8220 6072 9036 6100
rect 9030 6060 9036 6072
rect 9088 6100 9094 6112
rect 9508 6100 9536 6199
rect 10410 6196 10416 6248
rect 10468 6196 10474 6248
rect 9677 6171 9735 6177
rect 9677 6137 9689 6171
rect 9723 6168 9735 6171
rect 11072 6168 11100 6267
rect 9723 6140 11100 6168
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 10502 6100 10508 6112
rect 9088 6072 10508 6100
rect 9088 6060 9094 6072
rect 10502 6060 10508 6072
rect 10560 6100 10566 6112
rect 10689 6103 10747 6109
rect 10689 6100 10701 6103
rect 10560 6072 10701 6100
rect 10560 6060 10566 6072
rect 10689 6069 10701 6072
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 10778 6060 10784 6112
rect 10836 6100 10842 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10836 6072 10885 6100
rect 10836 6060 10842 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 10873 6063 10931 6069
rect 1104 6010 18124 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 18124 6010
rect 1104 5936 18124 5958
rect 2130 5856 2136 5908
rect 2188 5856 2194 5908
rect 2593 5899 2651 5905
rect 2593 5865 2605 5899
rect 2639 5896 2651 5899
rect 4062 5896 4068 5908
rect 2639 5868 4068 5896
rect 2639 5865 2651 5868
rect 2593 5859 2651 5865
rect 2608 5828 2636 5859
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4798 5896 4804 5908
rect 4448 5868 4804 5896
rect 3510 5828 3516 5840
rect 1872 5800 2636 5828
rect 2746 5800 3516 5828
rect 1872 5701 1900 5800
rect 2746 5760 2774 5800
rect 3510 5788 3516 5800
rect 3568 5788 3574 5840
rect 2516 5732 2774 5760
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 1946 5652 1952 5704
rect 2004 5652 2010 5704
rect 2516 5701 2544 5732
rect 2958 5720 2964 5772
rect 3016 5720 3022 5772
rect 3050 5720 3056 5772
rect 3108 5720 3114 5772
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5760 3295 5763
rect 3694 5760 3700 5772
rect 3283 5732 3700 5760
rect 3283 5729 3295 5732
rect 3237 5723 3295 5729
rect 3694 5720 3700 5732
rect 3752 5720 3758 5772
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 4028 5732 4292 5760
rect 4028 5720 4034 5732
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 2056 5664 2329 5692
rect 1670 5584 1676 5636
rect 1728 5624 1734 5636
rect 2056 5624 2084 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 2516 5695 2578 5701
rect 2516 5664 2532 5695
rect 2317 5655 2375 5661
rect 2520 5661 2532 5664
rect 2566 5661 2578 5695
rect 2520 5655 2578 5661
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5692 2743 5695
rect 2774 5692 2780 5704
rect 2731 5664 2780 5692
rect 2731 5661 2743 5664
rect 2685 5655 2743 5661
rect 2774 5652 2780 5664
rect 2832 5692 2838 5704
rect 3145 5695 3203 5701
rect 2832 5664 2912 5692
rect 2832 5652 2838 5664
rect 1728 5596 2084 5624
rect 2133 5627 2191 5633
rect 1728 5584 1734 5596
rect 2133 5593 2145 5627
rect 2179 5624 2191 5627
rect 2884 5624 2912 5664
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 3160 5624 3188 5655
rect 3510 5652 3516 5704
rect 3568 5692 3574 5704
rect 4264 5701 4292 5732
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 3568 5664 4169 5692
rect 3568 5652 3574 5664
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 4448 5692 4476 5868
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 13633 5899 13691 5905
rect 13633 5896 13645 5899
rect 12032 5868 13645 5896
rect 12032 5856 12038 5868
rect 13633 5865 13645 5868
rect 13679 5865 13691 5899
rect 13633 5859 13691 5865
rect 7745 5831 7803 5837
rect 7745 5797 7757 5831
rect 7791 5828 7803 5831
rect 11885 5831 11943 5837
rect 7791 5800 8432 5828
rect 7791 5797 7803 5800
rect 7745 5791 7803 5797
rect 6012 5732 6408 5760
rect 4387 5664 4476 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4614 5652 4620 5704
rect 4672 5692 4678 5704
rect 6012 5692 6040 5732
rect 4672 5664 6040 5692
rect 6089 5695 6147 5701
rect 4672 5652 4678 5664
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 3694 5624 3700 5636
rect 2179 5596 2820 5624
rect 2884 5596 3700 5624
rect 2179 5593 2191 5596
rect 2133 5587 2191 5593
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 2682 5556 2688 5568
rect 2455 5528 2688 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 2792 5565 2820 5596
rect 3694 5584 3700 5596
rect 3752 5584 3758 5636
rect 4525 5627 4583 5633
rect 4525 5593 4537 5627
rect 4571 5593 4583 5627
rect 4525 5587 4583 5593
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5525 2835 5559
rect 2777 5519 2835 5525
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5556 4031 5559
rect 4430 5556 4436 5568
rect 4019 5528 4436 5556
rect 4019 5525 4031 5528
rect 3973 5519 4031 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 4540 5556 4568 5587
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 4862 5627 4920 5633
rect 4862 5624 4874 5627
rect 4764 5596 4874 5624
rect 4764 5584 4770 5596
rect 4862 5593 4874 5596
rect 4908 5593 4920 5627
rect 4862 5587 4920 5593
rect 5534 5556 5540 5568
rect 4540 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5556 5598 5568
rect 5997 5559 6055 5565
rect 5997 5556 6009 5559
rect 5592 5528 6009 5556
rect 5592 5516 5598 5528
rect 5997 5525 6009 5528
rect 6043 5525 6055 5559
rect 6104 5556 6132 5655
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 6380 5701 6408 5732
rect 8404 5704 8432 5800
rect 11885 5797 11897 5831
rect 11931 5797 11943 5831
rect 11885 5791 11943 5797
rect 11701 5763 11759 5769
rect 11701 5760 11713 5763
rect 10980 5732 11713 5760
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6914 5692 6920 5704
rect 6411 5664 6920 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 6914 5652 6920 5664
rect 6972 5692 6978 5704
rect 7374 5692 7380 5704
rect 6972 5664 7380 5692
rect 6972 5652 6978 5664
rect 7374 5652 7380 5664
rect 7432 5652 7438 5704
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5692 9183 5695
rect 9306 5692 9312 5704
rect 9171 5664 9312 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 9398 5652 9404 5704
rect 9456 5652 9462 5704
rect 10778 5652 10784 5704
rect 10836 5701 10842 5704
rect 10836 5692 10848 5701
rect 10836 5664 10881 5692
rect 10836 5655 10848 5664
rect 10836 5652 10842 5655
rect 6181 5627 6239 5633
rect 6181 5593 6193 5627
rect 6227 5624 6239 5627
rect 6610 5627 6668 5633
rect 6610 5624 6622 5627
rect 6227 5596 6622 5624
rect 6227 5593 6239 5596
rect 6181 5587 6239 5593
rect 6610 5593 6622 5596
rect 6656 5593 6668 5627
rect 6610 5587 6668 5593
rect 7282 5584 7288 5636
rect 7340 5624 7346 5636
rect 7837 5627 7895 5633
rect 7837 5624 7849 5627
rect 7340 5596 7849 5624
rect 7340 5584 7346 5596
rect 7837 5593 7849 5596
rect 7883 5593 7895 5627
rect 7837 5587 7895 5593
rect 9030 5584 9036 5636
rect 9088 5624 9094 5636
rect 9217 5627 9275 5633
rect 9217 5624 9229 5627
rect 9088 5596 9229 5624
rect 9088 5584 9094 5596
rect 9217 5593 9229 5596
rect 9263 5593 9275 5627
rect 9217 5587 9275 5593
rect 10502 5584 10508 5636
rect 10560 5624 10566 5636
rect 10980 5624 11008 5732
rect 11701 5729 11713 5732
rect 11747 5729 11759 5763
rect 11900 5760 11928 5791
rect 11900 5732 12020 5760
rect 11701 5723 11759 5729
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 10560 5596 11008 5624
rect 11072 5624 11100 5655
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11388 5664 11529 5692
rect 11388 5652 11394 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 11606 5652 11612 5704
rect 11664 5652 11670 5704
rect 11882 5652 11888 5704
rect 11940 5652 11946 5704
rect 11992 5701 12020 5732
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 12158 5652 12164 5704
rect 12216 5652 12222 5704
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 12342 5692 12348 5704
rect 12299 5664 12348 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 12268 5624 12296 5655
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 12498 5627 12556 5633
rect 12498 5624 12510 5627
rect 11072 5596 12296 5624
rect 12406 5596 12510 5624
rect 10560 5584 10566 5596
rect 7098 5556 7104 5568
rect 6104 5528 7104 5556
rect 5997 5519 6055 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 8665 5559 8723 5565
rect 8665 5556 8677 5559
rect 8352 5528 8677 5556
rect 8352 5516 8358 5528
rect 8665 5525 8677 5528
rect 8711 5525 8723 5559
rect 8665 5519 8723 5525
rect 9582 5516 9588 5568
rect 9640 5516 9646 5568
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 10410 5556 10416 5568
rect 9723 5528 10416 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 11330 5516 11336 5568
rect 11388 5556 11394 5568
rect 11882 5556 11888 5568
rect 11388 5528 11888 5556
rect 11388 5516 11394 5528
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12069 5559 12127 5565
rect 12069 5525 12081 5559
rect 12115 5556 12127 5559
rect 12406 5556 12434 5596
rect 12498 5593 12510 5596
rect 12544 5593 12556 5627
rect 12498 5587 12556 5593
rect 12115 5528 12434 5556
rect 12115 5525 12127 5528
rect 12069 5519 12127 5525
rect 1104 5466 18124 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 18124 5466
rect 1104 5392 18124 5414
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3605 5355 3663 5361
rect 3605 5352 3617 5355
rect 3108 5324 3617 5352
rect 3108 5312 3114 5324
rect 3605 5321 3617 5324
rect 3651 5321 3663 5355
rect 3605 5315 3663 5321
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 4706 5352 4712 5364
rect 4203 5324 4712 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6733 5355 6791 5361
rect 6733 5352 6745 5355
rect 6328 5324 6745 5352
rect 6328 5312 6334 5324
rect 6733 5321 6745 5324
rect 6779 5321 6791 5355
rect 6733 5315 6791 5321
rect 7009 5355 7067 5361
rect 7009 5321 7021 5355
rect 7055 5352 7067 5355
rect 8294 5352 8300 5364
rect 7055 5324 8300 5352
rect 7055 5321 7067 5324
rect 7009 5315 7067 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 8389 5355 8447 5361
rect 8389 5321 8401 5355
rect 8435 5321 8447 5355
rect 8389 5315 8447 5321
rect 8665 5355 8723 5361
rect 8665 5321 8677 5355
rect 8711 5352 8723 5355
rect 8754 5352 8760 5364
rect 8711 5324 8760 5352
rect 8711 5321 8723 5324
rect 8665 5315 8723 5321
rect 4985 5287 5043 5293
rect 4985 5284 4997 5287
rect 3896 5256 4997 5284
rect 2958 5176 2964 5228
rect 3016 5216 3022 5228
rect 3513 5219 3571 5225
rect 3513 5216 3525 5219
rect 3016 5188 3525 5216
rect 3016 5176 3022 5188
rect 3513 5185 3525 5188
rect 3559 5216 3571 5219
rect 3786 5216 3792 5228
rect 3559 5188 3792 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 3896 5225 3924 5256
rect 4985 5253 4997 5256
rect 5031 5253 5043 5287
rect 4985 5247 5043 5253
rect 7190 5244 7196 5296
rect 7248 5244 7254 5296
rect 7558 5244 7564 5296
rect 7616 5244 7622 5296
rect 7745 5287 7803 5293
rect 7745 5284 7757 5287
rect 7668 5256 7757 5284
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 4295 5188 4384 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 3694 5108 3700 5160
rect 3752 5108 3758 5160
rect 4080 5148 4108 5179
rect 4356 5157 4384 5188
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4617 5219 4675 5225
rect 4617 5216 4629 5219
rect 4488 5188 4629 5216
rect 4488 5176 4494 5188
rect 4617 5185 4629 5188
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 5810 5216 5816 5228
rect 4847 5188 5816 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 5902 5176 5908 5228
rect 5960 5216 5966 5228
rect 6638 5216 6644 5228
rect 5960 5188 6644 5216
rect 5960 5176 5966 5188
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 6917 5219 6975 5225
rect 6917 5216 6929 5219
rect 6871 5188 6929 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 6917 5185 6929 5188
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 3896 5120 4108 5148
rect 4341 5151 4399 5157
rect 3712 5012 3740 5108
rect 3896 5089 3924 5120
rect 4341 5117 4353 5151
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5117 4583 5151
rect 4525 5111 4583 5117
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5117 4767 5151
rect 4709 5111 4767 5117
rect 3881 5083 3939 5089
rect 3881 5049 3893 5083
rect 3927 5049 3939 5083
rect 3881 5043 3939 5049
rect 3970 5040 3976 5092
rect 4028 5080 4034 5092
rect 4540 5080 4568 5111
rect 4028 5052 4568 5080
rect 4028 5040 4034 5052
rect 4062 5012 4068 5024
rect 3712 4984 4068 5012
rect 4062 4972 4068 4984
rect 4120 5012 4126 5024
rect 4724 5012 4752 5111
rect 5534 5108 5540 5160
rect 5592 5108 5598 5160
rect 4798 5040 4804 5092
rect 4856 5080 4862 5092
rect 5920 5080 5948 5176
rect 6932 5148 6960 5179
rect 7282 5176 7288 5228
rect 7340 5176 7346 5228
rect 7668 5225 7696 5256
rect 7745 5253 7757 5256
rect 7791 5284 7803 5287
rect 7791 5256 8248 5284
rect 7791 5253 7803 5256
rect 7745 5247 7803 5253
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 8110 5176 8116 5228
rect 8168 5176 8174 5228
rect 8220 5225 8248 5256
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 8294 5176 8300 5228
rect 8352 5176 8358 5228
rect 6932 5120 7420 5148
rect 4856 5052 5948 5080
rect 4856 5040 4862 5052
rect 7098 5040 7104 5092
rect 7156 5080 7162 5092
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 7156 5052 7297 5080
rect 7156 5040 7162 5052
rect 7285 5049 7297 5052
rect 7331 5049 7343 5083
rect 7392 5080 7420 5120
rect 7466 5108 7472 5160
rect 7524 5108 7530 5160
rect 8297 5083 8355 5089
rect 8297 5080 8309 5083
rect 7392 5052 8309 5080
rect 7285 5043 7343 5049
rect 8297 5049 8309 5052
rect 8343 5049 8355 5083
rect 8297 5043 8355 5049
rect 4120 4984 4752 5012
rect 4120 4972 4126 4984
rect 7190 4972 7196 5024
rect 7248 4972 7254 5024
rect 7558 4972 7564 5024
rect 7616 5012 7622 5024
rect 8404 5012 8432 5315
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 12158 5312 12164 5364
rect 12216 5352 12222 5364
rect 12253 5355 12311 5361
rect 12253 5352 12265 5355
rect 12216 5324 12265 5352
rect 12216 5312 12222 5324
rect 12253 5321 12265 5324
rect 12299 5321 12311 5355
rect 12253 5315 12311 5321
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5216 8631 5219
rect 9030 5216 9036 5228
rect 8619 5188 9036 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 9030 5176 9036 5188
rect 9088 5216 9094 5228
rect 9306 5216 9312 5228
rect 9088 5188 9312 5216
rect 9088 5176 9094 5188
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 12250 5176 12256 5228
rect 12308 5176 12314 5228
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5216 12495 5219
rect 12618 5216 12624 5228
rect 12483 5188 12624 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 8754 5108 8760 5160
rect 8812 5148 8818 5160
rect 9122 5148 9128 5160
rect 8812 5120 9128 5148
rect 8812 5108 8818 5120
rect 9122 5108 9128 5120
rect 9180 5148 9186 5160
rect 9217 5151 9275 5157
rect 9217 5148 9229 5151
rect 9180 5120 9229 5148
rect 9180 5108 9186 5120
rect 9217 5117 9229 5120
rect 9263 5117 9275 5151
rect 9217 5111 9275 5117
rect 7616 4984 8432 5012
rect 7616 4972 7622 4984
rect 1104 4922 18124 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 18124 4922
rect 1104 4848 18124 4870
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 13357 4811 13415 4817
rect 13357 4808 13369 4811
rect 12676 4780 13369 4808
rect 12676 4768 12682 4780
rect 13357 4777 13369 4780
rect 13403 4777 13415 4811
rect 13357 4771 13415 4777
rect 12802 4700 12808 4752
rect 12860 4700 12866 4752
rect 7190 4632 7196 4684
rect 7248 4672 7254 4684
rect 9217 4675 9275 4681
rect 7248 4644 7512 4672
rect 7248 4632 7254 4644
rect 7374 4564 7380 4616
rect 7432 4564 7438 4616
rect 7484 4604 7512 4644
rect 9217 4641 9229 4675
rect 9263 4672 9275 4675
rect 10042 4672 10048 4684
rect 9263 4644 10048 4672
rect 9263 4641 9275 4644
rect 9217 4635 9275 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 12492 4644 13216 4672
rect 12492 4632 12498 4644
rect 7633 4607 7691 4613
rect 7633 4604 7645 4607
rect 7484 4576 7645 4604
rect 7633 4573 7645 4576
rect 7679 4573 7691 4607
rect 7633 4567 7691 4573
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9140 4536 9168 4567
rect 9306 4564 9312 4616
rect 9364 4564 9370 4616
rect 9398 4564 9404 4616
rect 9456 4564 9462 4616
rect 12250 4564 12256 4616
rect 12308 4604 12314 4616
rect 13188 4613 13216 4644
rect 13081 4607 13139 4613
rect 13081 4604 13093 4607
rect 12308 4576 13093 4604
rect 12308 4564 12314 4576
rect 13081 4573 13093 4576
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4604 13231 4607
rect 13630 4604 13636 4616
rect 13219 4576 13636 4604
rect 13219 4573 13231 4576
rect 13173 4567 13231 4573
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 17770 4564 17776 4616
rect 17828 4564 17834 4616
rect 9950 4536 9956 4548
rect 9140 4508 9956 4536
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 12621 4539 12679 4545
rect 12621 4505 12633 4539
rect 12667 4505 12679 4539
rect 12621 4499 12679 4505
rect 3970 4428 3976 4480
rect 4028 4468 4034 4480
rect 6086 4468 6092 4480
rect 4028 4440 6092 4468
rect 4028 4428 4034 4440
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 8754 4428 8760 4480
rect 8812 4428 8818 4480
rect 8938 4428 8944 4480
rect 8996 4428 9002 4480
rect 12636 4468 12664 4499
rect 12710 4496 12716 4548
rect 12768 4536 12774 4548
rect 12805 4539 12863 4545
rect 12805 4536 12817 4539
rect 12768 4508 12817 4536
rect 12768 4496 12774 4508
rect 12805 4505 12817 4508
rect 12851 4505 12863 4539
rect 12805 4499 12863 4505
rect 12912 4508 17632 4536
rect 12912 4468 12940 4508
rect 12636 4440 12940 4468
rect 12986 4428 12992 4480
rect 13044 4428 13050 4480
rect 17604 4477 17632 4508
rect 17589 4471 17647 4477
rect 17589 4437 17601 4471
rect 17635 4437 17647 4471
rect 17589 4431 17647 4437
rect 1104 4378 18124 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 18124 4378
rect 1104 4304 18124 4326
rect 4249 4267 4307 4273
rect 4249 4233 4261 4267
rect 4295 4264 4307 4267
rect 4614 4264 4620 4276
rect 4295 4236 4620 4264
rect 4295 4233 4307 4236
rect 4249 4227 4307 4233
rect 4614 4224 4620 4236
rect 4672 4264 4678 4276
rect 5905 4267 5963 4273
rect 5905 4264 5917 4267
rect 4672 4236 5917 4264
rect 4672 4224 4678 4236
rect 5905 4233 5917 4236
rect 5951 4264 5963 4267
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 5951 4236 6561 4264
rect 5951 4233 5963 4236
rect 5905 4227 5963 4233
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 6638 4224 6644 4276
rect 6696 4264 6702 4276
rect 6917 4267 6975 4273
rect 6917 4264 6929 4267
rect 6696 4236 6929 4264
rect 6696 4224 6702 4236
rect 6917 4233 6929 4236
rect 6963 4233 6975 4267
rect 6917 4227 6975 4233
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 6932 4196 6960 4227
rect 10042 4224 10048 4276
rect 10100 4224 10106 4276
rect 10137 4267 10195 4273
rect 10137 4233 10149 4267
rect 10183 4264 10195 4267
rect 10778 4264 10784 4276
rect 10183 4236 10784 4264
rect 10183 4233 10195 4236
rect 10137 4227 10195 4233
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 11701 4267 11759 4273
rect 11701 4233 11713 4267
rect 11747 4264 11759 4267
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11747 4236 11989 4264
rect 11747 4233 11759 4236
rect 11701 4227 11759 4233
rect 11977 4233 11989 4236
rect 12023 4233 12035 4267
rect 11977 4227 12035 4233
rect 8113 4199 8171 4205
rect 4120 4168 5488 4196
rect 6932 4168 7328 4196
rect 4120 4156 4126 4168
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 4028 4100 4169 4128
rect 4028 4088 4034 4100
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 4356 4069 4384 4168
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 4709 4131 4767 4137
rect 4709 4097 4721 4131
rect 4755 4128 4767 4131
rect 4798 4128 4804 4140
rect 4755 4100 4804 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4540 4060 4568 4091
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 4893 4131 4951 4137
rect 4893 4097 4905 4131
rect 4939 4128 4951 4131
rect 4939 4100 5396 4128
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 4985 4063 5043 4069
rect 4985 4060 4997 4063
rect 4540 4032 4997 4060
rect 4341 4023 4399 4029
rect 4985 4029 4997 4032
rect 5031 4029 5043 4063
rect 4985 4023 5043 4029
rect 5368 3936 5396 4100
rect 5460 4060 5488 4168
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4128 5687 4131
rect 5902 4128 5908 4140
rect 5675 4100 5908 4128
rect 5675 4097 5687 4100
rect 5629 4091 5687 4097
rect 5902 4088 5908 4100
rect 5960 4128 5966 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5960 4100 6009 4128
rect 5960 4088 5966 4100
rect 5997 4097 6009 4100
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 6086 4088 6092 4140
rect 6144 4128 6150 4140
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 6144 4100 6653 4128
rect 6144 4088 6150 4100
rect 6641 4097 6653 4100
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 6730 4088 6736 4140
rect 6788 4088 6794 4140
rect 7098 4088 7104 4140
rect 7156 4088 7162 4140
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7300 4128 7328 4168
rect 8113 4165 8125 4199
rect 8159 4196 8171 4199
rect 8938 4196 8944 4208
rect 8159 4168 8944 4196
rect 8159 4165 8171 4168
rect 8113 4159 8171 4165
rect 8938 4156 8944 4168
rect 8996 4156 9002 4208
rect 10069 4196 10097 4224
rect 11606 4196 11612 4208
rect 10069 4168 11612 4196
rect 11606 4156 11612 4168
rect 11664 4196 11670 4208
rect 12802 4205 12808 4208
rect 11793 4199 11851 4205
rect 11793 4196 11805 4199
rect 11664 4168 11805 4196
rect 11664 4156 11670 4168
rect 11793 4165 11805 4168
rect 11839 4165 11851 4199
rect 12796 4196 12808 4205
rect 12763 4168 12808 4196
rect 11793 4159 11851 4165
rect 12796 4159 12808 4168
rect 12802 4156 12808 4159
rect 12860 4156 12866 4208
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 7300 4100 7389 4128
rect 7193 4091 7251 4097
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4128 7987 4131
rect 9030 4128 9036 4140
rect 7975 4100 9036 4128
rect 7975 4097 7987 4100
rect 7929 4091 7987 4097
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 5460 4032 5733 4060
rect 5721 4029 5733 4032
rect 5767 4060 5779 4063
rect 6365 4063 6423 4069
rect 6365 4060 6377 4063
rect 5767 4032 6377 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6365 4029 6377 4032
rect 6411 4029 6423 4063
rect 6365 4023 6423 4029
rect 7006 4020 7012 4072
rect 7064 4060 7070 4072
rect 7208 4060 7236 4091
rect 7852 4060 7880 4091
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 10244 4100 11744 4128
rect 10244 4060 10272 4100
rect 7064 4032 7880 4060
rect 8036 4032 10272 4060
rect 10321 4063 10379 4069
rect 7064 4020 7070 4032
rect 7282 3952 7288 4004
rect 7340 3952 7346 4004
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 4614 3924 4620 3936
rect 4571 3896 4620 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4798 3884 4804 3936
rect 4856 3884 4862 3936
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 5813 3927 5871 3933
rect 5813 3924 5825 3927
rect 5408 3896 5825 3924
rect 5408 3884 5414 3896
rect 5813 3893 5825 3896
rect 5859 3893 5871 3927
rect 5813 3887 5871 3893
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 7006 3924 7012 3936
rect 6687 3896 7012 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 8036 3924 8064 4032
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 10502 4060 10508 4072
rect 10367 4032 10508 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 11054 4020 11060 4072
rect 11112 4020 11118 4072
rect 11517 4063 11575 4069
rect 11517 4029 11529 4063
rect 11563 4029 11575 4063
rect 11716 4060 11744 4100
rect 11882 4088 11888 4140
rect 11940 4088 11946 4140
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 12032 4100 12173 4128
rect 12032 4088 12038 4100
rect 12161 4097 12173 4100
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4128 12403 4131
rect 12391 4100 12480 4128
rect 12391 4097 12403 4100
rect 12345 4091 12403 4097
rect 12452 4072 12480 4100
rect 12526 4088 12532 4140
rect 12584 4088 12590 4140
rect 12636 4100 13952 4128
rect 12250 4060 12256 4072
rect 11716 4032 12256 4060
rect 11517 4023 11575 4029
rect 10045 3995 10103 4001
rect 10045 3961 10057 3995
rect 10091 3992 10103 3995
rect 11238 3992 11244 4004
rect 10091 3964 11244 3992
rect 10091 3961 10103 3964
rect 10045 3955 10103 3961
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 7156 3896 8064 3924
rect 7156 3884 7162 3896
rect 8110 3884 8116 3936
rect 8168 3884 8174 3936
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 10284 3896 10425 3924
rect 10284 3884 10290 3896
rect 10413 3893 10425 3896
rect 10459 3893 10471 3927
rect 10413 3887 10471 3893
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 11532 3924 11560 4023
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 12636 4060 12664 4100
rect 12492 4032 12664 4060
rect 13924 4060 13952 4100
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 13924 4032 14565 4060
rect 12492 4020 12498 4032
rect 13924 4001 13952 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 13909 3995 13967 4001
rect 13909 3961 13921 3995
rect 13955 3961 13967 3995
rect 13909 3955 13967 3961
rect 10560 3896 11560 3924
rect 11793 3927 11851 3933
rect 10560 3884 10566 3896
rect 11793 3893 11805 3927
rect 11839 3924 11851 3927
rect 12342 3924 12348 3936
rect 11839 3896 12348 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 13998 3884 14004 3936
rect 14056 3884 14062 3936
rect 1104 3834 18124 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 18124 3834
rect 1104 3760 18124 3782
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 6788 3692 7941 3720
rect 6788 3680 6794 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 9030 3680 9036 3732
rect 9088 3680 9094 3732
rect 10318 3680 10324 3732
rect 10376 3720 10382 3732
rect 10597 3723 10655 3729
rect 10597 3720 10609 3723
rect 10376 3692 10609 3720
rect 10376 3680 10382 3692
rect 10597 3689 10609 3692
rect 10643 3689 10655 3723
rect 10597 3683 10655 3689
rect 12529 3723 12587 3729
rect 12529 3689 12541 3723
rect 12575 3720 12587 3723
rect 12710 3720 12716 3732
rect 12575 3692 12716 3720
rect 12575 3689 12587 3692
rect 12529 3683 12587 3689
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 12805 3723 12863 3729
rect 12805 3689 12817 3723
rect 12851 3720 12863 3723
rect 12986 3720 12992 3732
rect 12851 3692 12992 3720
rect 12851 3689 12863 3692
rect 12805 3683 12863 3689
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 4614 3612 4620 3664
rect 4672 3612 4678 3664
rect 5629 3655 5687 3661
rect 5629 3621 5641 3655
rect 5675 3652 5687 3655
rect 5718 3652 5724 3664
rect 5675 3624 5724 3652
rect 5675 3621 5687 3624
rect 5629 3615 5687 3621
rect 5718 3612 5724 3624
rect 5776 3612 5782 3664
rect 9490 3612 9496 3664
rect 9548 3612 9554 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 11882 3652 11888 3664
rect 10008 3624 11888 3652
rect 10008 3612 10014 3624
rect 11882 3612 11888 3624
rect 11940 3612 11946 3664
rect 12434 3652 12440 3664
rect 12406 3612 12440 3652
rect 12492 3612 12498 3664
rect 4632 3584 4660 3612
rect 4448 3556 4660 3584
rect 4448 3525 4476 3556
rect 7926 3544 7932 3596
rect 7984 3584 7990 3596
rect 11238 3584 11244 3596
rect 7984 3556 8800 3584
rect 7984 3544 7990 3556
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 4798 3516 4804 3528
rect 4663 3488 4804 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5350 3476 5356 3528
rect 5408 3476 5414 3528
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 5828 3516 5948 3518
rect 7374 3516 7380 3528
rect 5776 3490 7380 3516
rect 5776 3488 5856 3490
rect 5920 3488 7380 3490
rect 5776 3476 5782 3488
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 5810 3408 5816 3460
rect 5868 3448 5874 3460
rect 5966 3451 6024 3457
rect 5966 3448 5978 3451
rect 5868 3420 5978 3448
rect 5868 3408 5874 3420
rect 5966 3417 5978 3420
rect 6012 3417 6024 3451
rect 7760 3448 7788 3479
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 8772 3525 8800 3556
rect 9784 3556 11244 3584
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 7892 3488 8125 3516
rect 7892 3476 7898 3488
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 8220 3448 8248 3479
rect 9122 3476 9128 3528
rect 9180 3476 9186 3528
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3516 9551 3519
rect 9582 3516 9588 3528
rect 9539 3488 9588 3516
rect 9539 3485 9551 3488
rect 9493 3479 9551 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9784 3525 9812 3556
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 12406 3584 12434 3612
rect 11532 3556 12434 3584
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 10226 3476 10232 3528
rect 10284 3476 10290 3528
rect 10689 3519 10747 3525
rect 10689 3485 10701 3519
rect 10735 3516 10747 3519
rect 10735 3488 10916 3516
rect 10735 3485 10747 3488
rect 10689 3479 10747 3485
rect 5966 3411 6024 3417
rect 7116 3420 8248 3448
rect 10888 3448 10916 3488
rect 11146 3476 11152 3528
rect 11204 3476 11210 3528
rect 11532 3525 11560 3556
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3485 11575 3519
rect 11517 3479 11575 3485
rect 11882 3476 11888 3528
rect 11940 3476 11946 3528
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12437 3519 12495 3525
rect 12437 3516 12449 3519
rect 12400 3488 12449 3516
rect 12400 3476 12406 3488
rect 12437 3485 12449 3488
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 12618 3476 12624 3528
rect 12676 3476 12682 3528
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 13998 3516 14004 3528
rect 12943 3488 14004 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 11054 3448 11060 3460
rect 10888 3420 11060 3448
rect 4522 3340 4528 3392
rect 4580 3340 4586 3392
rect 5445 3383 5503 3389
rect 5445 3349 5457 3383
rect 5491 3380 5503 3383
rect 6454 3380 6460 3392
rect 5491 3352 6460 3380
rect 5491 3349 5503 3352
rect 5445 3343 5503 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7116 3389 7144 3420
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 11606 3408 11612 3460
rect 11664 3448 11670 3460
rect 12069 3451 12127 3457
rect 12069 3448 12081 3451
rect 11664 3420 12081 3448
rect 11664 3408 11670 3420
rect 12069 3417 12081 3420
rect 12115 3417 12127 3451
rect 12069 3411 12127 3417
rect 7101 3383 7159 3389
rect 7101 3380 7113 3383
rect 6972 3352 7113 3380
rect 6972 3340 6978 3352
rect 7101 3349 7113 3352
rect 7147 3349 7159 3383
rect 7101 3343 7159 3349
rect 7190 3340 7196 3392
rect 7248 3340 7254 3392
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 8573 3383 8631 3389
rect 8573 3380 8585 3383
rect 8444 3352 8585 3380
rect 8444 3340 8450 3352
rect 8573 3349 8585 3352
rect 8619 3349 8631 3383
rect 8573 3343 8631 3349
rect 9677 3383 9735 3389
rect 9677 3349 9689 3383
rect 9723 3380 9735 3383
rect 10137 3383 10195 3389
rect 10137 3380 10149 3383
rect 9723 3352 10149 3380
rect 9723 3349 9735 3352
rect 9677 3343 9735 3349
rect 10137 3349 10149 3352
rect 10183 3349 10195 3383
rect 10137 3343 10195 3349
rect 12158 3340 12164 3392
rect 12216 3389 12222 3392
rect 12216 3343 12225 3389
rect 12253 3383 12311 3389
rect 12253 3349 12265 3383
rect 12299 3380 12311 3383
rect 13538 3380 13544 3392
rect 12299 3352 13544 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 12216 3340 12222 3343
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 1104 3290 18124 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 18124 3290
rect 1104 3216 18124 3238
rect 6454 3136 6460 3188
rect 6512 3136 6518 3188
rect 9122 3136 9128 3188
rect 9180 3136 9186 3188
rect 10597 3179 10655 3185
rect 10597 3145 10609 3179
rect 10643 3176 10655 3179
rect 11054 3176 11060 3188
rect 10643 3148 11060 3176
rect 10643 3145 10655 3148
rect 10597 3139 10655 3145
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 11606 3136 11612 3188
rect 11664 3136 11670 3188
rect 12618 3176 12624 3188
rect 11716 3148 12624 3176
rect 4148 3111 4206 3117
rect 4148 3077 4160 3111
rect 4194 3108 4206 3111
rect 4522 3108 4528 3120
rect 4194 3080 4528 3108
rect 4194 3077 4206 3080
rect 4148 3071 4206 3077
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 7190 3108 7196 3120
rect 6564 3080 7196 3108
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 5718 3040 5724 3052
rect 3927 3012 5724 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 6564 3049 6592 3080
rect 7190 3068 7196 3080
rect 7248 3068 7254 3120
rect 7834 3108 7840 3120
rect 7392 3080 7840 3108
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 5534 2932 5540 2984
rect 5592 2972 5598 2984
rect 6748 2972 6776 3003
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 7392 3049 7420 3080
rect 7834 3068 7840 3080
rect 7892 3068 7898 3120
rect 9490 3117 9496 3120
rect 9484 3108 9496 3117
rect 9451 3080 9496 3108
rect 9484 3071 9496 3080
rect 9490 3068 9496 3071
rect 9548 3068 9554 3120
rect 10949 3111 11007 3117
rect 10949 3077 10961 3111
rect 10995 3108 11007 3111
rect 10995 3080 11100 3108
rect 10995 3077 11007 3080
rect 10949 3071 11007 3077
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 6880 3012 7389 3040
rect 6880 3000 6886 3012
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 5592 2944 6776 2972
rect 5592 2932 5598 2944
rect 6914 2932 6920 2984
rect 6972 2972 6978 2984
rect 7484 2972 7512 3003
rect 6972 2944 7512 2972
rect 8220 2972 8248 3003
rect 8570 2972 8576 2984
rect 8220 2944 8576 2972
rect 6972 2932 6978 2944
rect 8570 2932 8576 2944
rect 8628 2932 8634 2984
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2941 9275 2975
rect 11072 2972 11100 3080
rect 11146 3068 11152 3120
rect 11204 3068 11210 3120
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11716 3049 11744 3148
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 12584 3080 13216 3108
rect 12584 3068 12590 3080
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11296 3012 11529 3040
rect 11296 3000 11302 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 12158 3000 12164 3052
rect 12216 3040 12222 3052
rect 13188 3049 13216 3080
rect 12906 3043 12964 3049
rect 12906 3040 12918 3043
rect 12216 3012 12918 3040
rect 12216 3000 12222 3012
rect 12906 3009 12918 3012
rect 12952 3009 12964 3043
rect 12906 3003 12964 3009
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 11882 2972 11888 2984
rect 11072 2944 11888 2972
rect 9217 2935 9275 2941
rect 7374 2864 7380 2916
rect 7432 2904 7438 2916
rect 9232 2904 9260 2935
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 7432 2876 9260 2904
rect 7432 2864 7438 2876
rect 10778 2864 10784 2916
rect 10836 2864 10842 2916
rect 10980 2876 11928 2904
rect 5261 2839 5319 2845
rect 5261 2805 5273 2839
rect 5307 2836 5319 2839
rect 5902 2836 5908 2848
rect 5307 2808 5908 2836
rect 5307 2805 5319 2808
rect 5261 2799 5319 2805
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 8113 2839 8171 2845
rect 8113 2805 8125 2839
rect 8159 2836 8171 2839
rect 9398 2836 9404 2848
rect 8159 2808 9404 2836
rect 8159 2805 8171 2808
rect 8113 2799 8171 2805
rect 9398 2796 9404 2808
rect 9456 2796 9462 2848
rect 10980 2845 11008 2876
rect 10965 2839 11023 2845
rect 10965 2805 10977 2839
rect 11011 2805 11023 2839
rect 10965 2799 11023 2805
rect 11146 2796 11152 2848
rect 11204 2836 11210 2848
rect 11790 2836 11796 2848
rect 11204 2808 11796 2836
rect 11204 2796 11210 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 11900 2836 11928 2876
rect 12434 2836 12440 2848
rect 11900 2808 12440 2836
rect 12434 2796 12440 2808
rect 12492 2836 12498 2848
rect 13354 2836 13360 2848
rect 12492 2808 13360 2836
rect 12492 2796 12498 2808
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 1104 2746 18124 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 18124 2746
rect 1104 2672 18124 2694
rect 13538 2592 13544 2644
rect 13596 2592 13602 2644
rect 8570 2524 8576 2576
rect 8628 2564 8634 2576
rect 8757 2567 8815 2573
rect 8757 2564 8769 2567
rect 8628 2536 8769 2564
rect 8628 2524 8634 2536
rect 8757 2533 8769 2536
rect 8803 2564 8815 2567
rect 8803 2536 9812 2564
rect 8803 2533 8815 2536
rect 8757 2527 8815 2533
rect 7374 2456 7380 2508
rect 7432 2456 7438 2508
rect 5534 2388 5540 2440
rect 5592 2388 5598 2440
rect 5902 2388 5908 2440
rect 5960 2428 5966 2440
rect 6822 2428 6828 2440
rect 5960 2400 6828 2428
rect 5960 2388 5966 2400
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 6914 2388 6920 2440
rect 6972 2388 6978 2440
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 7644 2431 7702 2437
rect 7644 2397 7656 2431
rect 7690 2428 7702 2431
rect 8110 2428 8116 2440
rect 7690 2400 8116 2428
rect 7690 2397 7702 2400
rect 7644 2391 7702 2397
rect 7300 2360 7328 2391
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 9784 2437 9812 2536
rect 12250 2524 12256 2576
rect 12308 2564 12314 2576
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 12308 2536 12817 2564
rect 12308 2524 12314 2536
rect 12805 2533 12817 2536
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 12667 2468 13492 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8812 2400 9137 2428
rect 8812 2388 8818 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 10410 2388 10416 2440
rect 10468 2388 10474 2440
rect 11054 2388 11060 2440
rect 11112 2388 11118 2440
rect 11882 2388 11888 2440
rect 11940 2428 11946 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11940 2400 11989 2428
rect 11940 2388 11946 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12066 2388 12072 2440
rect 12124 2428 12130 2440
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12124 2400 13001 2428
rect 12124 2388 12130 2400
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13354 2388 13360 2440
rect 13412 2388 13418 2440
rect 13464 2437 13492 2468
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 8294 2360 8300 2372
rect 7300 2332 8300 2360
rect 8294 2320 8300 2332
rect 8352 2320 8358 2372
rect 5721 2295 5779 2301
rect 5721 2261 5733 2295
rect 5767 2292 5779 2295
rect 5810 2292 5816 2304
rect 5767 2264 5816 2292
rect 5767 2261 5779 2264
rect 5721 2255 5779 2261
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 6089 2295 6147 2301
rect 6089 2261 6101 2295
rect 6135 2292 6147 2295
rect 6454 2292 6460 2304
rect 6135 2264 6460 2292
rect 6135 2261 6147 2264
rect 6089 2255 6147 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 6733 2295 6791 2301
rect 6733 2261 6745 2295
rect 6779 2292 6791 2295
rect 7006 2292 7012 2304
rect 6779 2264 7012 2292
rect 6779 2261 6791 2264
rect 6733 2255 6791 2261
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7101 2295 7159 2301
rect 7101 2261 7113 2295
rect 7147 2292 7159 2295
rect 7742 2292 7748 2304
rect 7147 2264 7748 2292
rect 7147 2261 7159 2264
rect 7101 2255 7159 2261
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 9732 2264 9965 2292
rect 9732 2252 9738 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 9953 2255 10011 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 10376 2264 10609 2292
rect 10376 2252 10382 2264
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 10597 2255 10655 2261
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 11241 2295 11299 2301
rect 11241 2292 11253 2295
rect 11020 2264 11253 2292
rect 11020 2252 11026 2264
rect 11241 2261 11253 2264
rect 11287 2261 11299 2295
rect 11241 2255 11299 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11664 2264 11713 2292
rect 11664 2252 11670 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 1104 2202 18124 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 18124 2202
rect 1104 2128 18124 2150
<< via1 >>
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 8576 18955 8628 18964
rect 8576 18921 8585 18955
rect 8585 18921 8619 18955
rect 8619 18921 8628 18955
rect 8576 18912 8628 18921
rect 9220 18955 9272 18964
rect 9220 18921 9229 18955
rect 9229 18921 9263 18955
rect 9263 18921 9272 18955
rect 9220 18912 9272 18921
rect 10876 18912 10928 18964
rect 11888 18955 11940 18964
rect 11888 18921 11897 18955
rect 11897 18921 11931 18955
rect 11931 18921 11940 18955
rect 11888 18912 11940 18921
rect 8760 18751 8812 18760
rect 8760 18717 8769 18751
rect 8769 18717 8803 18751
rect 8803 18717 8812 18751
rect 8760 18708 8812 18717
rect 9588 18708 9640 18760
rect 11336 18751 11388 18760
rect 11336 18717 11345 18751
rect 11345 18717 11379 18751
rect 11379 18717 11388 18751
rect 11336 18708 11388 18717
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 11336 14603 11388 14612
rect 11336 14569 11345 14603
rect 11345 14569 11379 14603
rect 11379 14569 11388 14603
rect 11336 14560 11388 14569
rect 848 14492 900 14544
rect 4804 14356 4856 14408
rect 6276 14356 6328 14408
rect 12900 14356 12952 14408
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 10232 14331 10284 14340
rect 10232 14297 10266 14331
rect 10266 14297 10284 14331
rect 10232 14288 10284 14297
rect 6736 14220 6788 14272
rect 14556 14220 14608 14272
rect 17684 14263 17736 14272
rect 17684 14229 17693 14263
rect 17693 14229 17727 14263
rect 17727 14229 17736 14263
rect 17684 14220 17736 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 2136 14016 2188 14068
rect 4804 14059 4856 14068
rect 4804 14025 4813 14059
rect 4813 14025 4847 14059
rect 4847 14025 4856 14059
rect 4804 14016 4856 14025
rect 8760 14059 8812 14068
rect 8760 14025 8769 14059
rect 8769 14025 8803 14059
rect 8803 14025 8812 14059
rect 8760 14016 8812 14025
rect 8944 14016 8996 14068
rect 11336 14016 11388 14068
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 7104 13948 7156 14000
rect 6736 13923 6788 13932
rect 6736 13889 6745 13923
rect 6745 13889 6779 13923
rect 6779 13889 6788 13923
rect 6736 13880 6788 13889
rect 8116 13880 8168 13932
rect 9128 13880 9180 13932
rect 11704 14016 11756 14068
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 10324 13923 10376 13932
rect 10324 13889 10333 13923
rect 10333 13889 10367 13923
rect 10367 13889 10376 13923
rect 10324 13880 10376 13889
rect 12624 13923 12676 13932
rect 12624 13889 12642 13923
rect 12642 13889 12676 13923
rect 12624 13880 12676 13889
rect 12900 13923 12952 13932
rect 12900 13889 12909 13923
rect 12909 13889 12943 13923
rect 12943 13889 12952 13923
rect 12900 13880 12952 13889
rect 13912 13880 13964 13932
rect 15200 13948 15252 14000
rect 15476 14016 15528 14068
rect 16120 14016 16172 14068
rect 17684 14059 17736 14068
rect 17684 14025 17693 14059
rect 17693 14025 17727 14059
rect 17727 14025 17736 14059
rect 17684 14016 17736 14025
rect 14924 13880 14976 13932
rect 6920 13812 6972 13864
rect 9312 13744 9364 13796
rect 11152 13744 11204 13796
rect 8852 13719 8904 13728
rect 8852 13685 8861 13719
rect 8861 13685 8895 13719
rect 8895 13685 8904 13719
rect 8852 13676 8904 13685
rect 9864 13719 9916 13728
rect 9864 13685 9873 13719
rect 9873 13685 9907 13719
rect 9907 13685 9916 13719
rect 9864 13676 9916 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 6368 13472 6420 13524
rect 10232 13472 10284 13524
rect 8944 13447 8996 13456
rect 8944 13413 8953 13447
rect 8953 13413 8987 13447
rect 8987 13413 8996 13447
rect 8944 13404 8996 13413
rect 12072 13404 12124 13456
rect 6552 13336 6604 13388
rect 7472 13336 7524 13388
rect 11704 13379 11756 13388
rect 11704 13345 11713 13379
rect 11713 13345 11747 13379
rect 11747 13345 11756 13379
rect 11704 13336 11756 13345
rect 12992 13472 13044 13524
rect 13912 13472 13964 13524
rect 14924 13472 14976 13524
rect 13636 13336 13688 13388
rect 4620 13268 4672 13320
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7012 13268 7064 13277
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 9496 13268 9548 13320
rect 9864 13311 9916 13320
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 11888 13268 11940 13320
rect 10508 13243 10560 13252
rect 10508 13209 10517 13243
rect 10517 13209 10551 13243
rect 10551 13209 10560 13243
rect 10508 13200 10560 13209
rect 13452 13243 13504 13252
rect 13452 13209 13461 13243
rect 13461 13209 13495 13243
rect 13495 13209 13504 13243
rect 14556 13311 14608 13320
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 14832 13311 14884 13320
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 15844 13268 15896 13320
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 13452 13200 13504 13209
rect 848 13132 900 13184
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 9404 13132 9456 13184
rect 10600 13132 10652 13184
rect 11704 13132 11756 13184
rect 14372 13132 14424 13184
rect 17316 13175 17368 13184
rect 17316 13141 17325 13175
rect 17325 13141 17359 13175
rect 17359 13141 17368 13175
rect 17316 13132 17368 13141
rect 17684 13175 17736 13184
rect 17684 13141 17693 13175
rect 17693 13141 17727 13175
rect 17727 13141 17736 13175
rect 17684 13132 17736 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 6368 12903 6420 12912
rect 6368 12869 6377 12903
rect 6377 12869 6411 12903
rect 6411 12869 6420 12903
rect 6368 12860 6420 12869
rect 5540 12792 5592 12844
rect 7104 12971 7156 12980
rect 7104 12937 7113 12971
rect 7113 12937 7147 12971
rect 7147 12937 7156 12971
rect 7104 12928 7156 12937
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 10508 12860 10560 12912
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 9312 12835 9364 12844
rect 9312 12801 9321 12835
rect 9321 12801 9355 12835
rect 9355 12801 9364 12835
rect 9312 12792 9364 12801
rect 11520 12860 11572 12912
rect 12072 12860 12124 12912
rect 13452 12928 13504 12980
rect 13268 12860 13320 12912
rect 11060 12835 11112 12844
rect 11060 12801 11069 12835
rect 11069 12801 11103 12835
rect 11103 12801 11112 12835
rect 11060 12792 11112 12801
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 14832 12792 14884 12844
rect 15936 12792 15988 12844
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 7748 12767 7800 12776
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 8852 12724 8904 12776
rect 10232 12724 10284 12776
rect 14740 12724 14792 12776
rect 17500 12767 17552 12776
rect 17500 12733 17509 12767
rect 17509 12733 17543 12767
rect 17543 12733 17552 12767
rect 17500 12724 17552 12733
rect 12624 12656 12676 12708
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 6644 12588 6696 12640
rect 7196 12588 7248 12640
rect 7748 12588 7800 12640
rect 10324 12588 10376 12640
rect 13820 12588 13872 12640
rect 16028 12631 16080 12640
rect 16028 12597 16037 12631
rect 16037 12597 16071 12631
rect 16071 12597 16080 12631
rect 16028 12588 16080 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 6368 12384 6420 12436
rect 8208 12384 8260 12436
rect 9036 12384 9088 12436
rect 14372 12427 14424 12436
rect 14372 12393 14381 12427
rect 14381 12393 14415 12427
rect 14415 12393 14424 12427
rect 14372 12384 14424 12393
rect 17500 12384 17552 12436
rect 6276 12359 6328 12368
rect 6276 12325 6285 12359
rect 6285 12325 6319 12359
rect 6319 12325 6328 12359
rect 6276 12316 6328 12325
rect 6552 12316 6604 12368
rect 4620 12180 4672 12232
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 7012 12248 7064 12300
rect 14832 12316 14884 12368
rect 7748 12248 7800 12300
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 6276 12180 6328 12232
rect 6368 12180 6420 12232
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 8392 12180 8444 12232
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 13268 12291 13320 12300
rect 13268 12257 13277 12291
rect 13277 12257 13311 12291
rect 13311 12257 13320 12291
rect 13268 12248 13320 12257
rect 14464 12248 14516 12300
rect 12808 12180 12860 12232
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 5632 12112 5684 12164
rect 8944 12112 8996 12164
rect 9588 12112 9640 12164
rect 12992 12155 13044 12164
rect 12992 12121 13001 12155
rect 13001 12121 13035 12155
rect 13035 12121 13044 12155
rect 12992 12112 13044 12121
rect 4620 12044 4672 12096
rect 5448 12044 5500 12096
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 6552 12044 6604 12053
rect 7012 12044 7064 12096
rect 8760 12044 8812 12096
rect 9220 12087 9272 12096
rect 9220 12053 9245 12087
rect 9245 12053 9272 12087
rect 9220 12044 9272 12053
rect 9404 12087 9456 12096
rect 9404 12053 9413 12087
rect 9413 12053 9447 12087
rect 9447 12053 9456 12087
rect 9404 12044 9456 12053
rect 11428 12044 11480 12096
rect 11612 12044 11664 12096
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15200 12248 15252 12300
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 15476 12112 15528 12164
rect 14740 12044 14792 12096
rect 15384 12044 15436 12096
rect 16212 12223 16264 12232
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 16028 12112 16080 12164
rect 17500 12044 17552 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 4712 11840 4764 11892
rect 6276 11840 6328 11892
rect 7656 11840 7708 11892
rect 8300 11840 8352 11892
rect 8760 11840 8812 11892
rect 9220 11840 9272 11892
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 10600 11883 10652 11892
rect 10600 11849 10609 11883
rect 10609 11849 10643 11883
rect 10643 11849 10652 11883
rect 10600 11840 10652 11849
rect 12808 11840 12860 11892
rect 15844 11840 15896 11892
rect 3884 11747 3936 11756
rect 3884 11713 3918 11747
rect 3918 11713 3936 11747
rect 3884 11704 3936 11713
rect 5448 11772 5500 11824
rect 5724 11772 5776 11824
rect 8392 11815 8444 11824
rect 8392 11781 8401 11815
rect 8401 11781 8435 11815
rect 8435 11781 8444 11815
rect 8392 11772 8444 11781
rect 8668 11772 8720 11824
rect 5632 11704 5684 11756
rect 6368 11704 6420 11756
rect 7012 11704 7064 11756
rect 8208 11704 8260 11756
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 8300 11568 8352 11620
rect 848 11500 900 11552
rect 9036 11704 9088 11756
rect 9404 11772 9456 11824
rect 9312 11704 9364 11756
rect 8668 11568 8720 11620
rect 9588 11704 9640 11756
rect 10048 11704 10100 11756
rect 11428 11772 11480 11824
rect 11244 11704 11296 11756
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 14832 11772 14884 11824
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12808 11747 12860 11756
rect 12808 11713 12817 11747
rect 12817 11713 12851 11747
rect 12851 11713 12860 11747
rect 12808 11704 12860 11713
rect 14924 11704 14976 11756
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 16120 11704 16172 11756
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 15384 11636 15436 11688
rect 17132 11679 17184 11688
rect 17132 11645 17141 11679
rect 17141 11645 17175 11679
rect 17175 11645 17184 11679
rect 17132 11636 17184 11645
rect 17776 11636 17828 11688
rect 10048 11568 10100 11620
rect 14556 11568 14608 11620
rect 9404 11500 9456 11552
rect 9772 11500 9824 11552
rect 12072 11500 12124 11552
rect 14832 11500 14884 11552
rect 16672 11543 16724 11552
rect 16672 11509 16681 11543
rect 16681 11509 16715 11543
rect 16715 11509 16724 11543
rect 16672 11500 16724 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 3884 11296 3936 11348
rect 4712 11296 4764 11348
rect 6460 11296 6512 11348
rect 7472 11296 7524 11348
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 14556 11296 14608 11348
rect 15936 11296 15988 11348
rect 17776 11339 17828 11348
rect 17776 11305 17785 11339
rect 17785 11305 17819 11339
rect 17819 11305 17828 11339
rect 17776 11296 17828 11305
rect 4620 11228 4672 11280
rect 9680 11228 9732 11280
rect 4528 11135 4580 11144
rect 4528 11101 4537 11135
rect 4537 11101 4571 11135
rect 4571 11101 4580 11135
rect 4528 11092 4580 11101
rect 4712 11092 4764 11144
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 6552 11092 6604 11144
rect 9220 11160 9272 11212
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9496 11160 9548 11212
rect 14372 11228 14424 11280
rect 16120 11228 16172 11280
rect 9404 11092 9456 11144
rect 6736 11024 6788 11076
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 11152 11092 11204 11144
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 12164 11092 12216 11144
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 15292 11160 15344 11212
rect 12624 11092 12676 11144
rect 13084 11092 13136 11144
rect 14924 11135 14976 11144
rect 14924 11101 14933 11135
rect 14933 11101 14967 11135
rect 14967 11101 14976 11135
rect 14924 11092 14976 11101
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 16212 11092 16264 11144
rect 16672 11135 16724 11144
rect 16672 11101 16706 11135
rect 16706 11101 16724 11135
rect 16672 11092 16724 11101
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 6828 10956 6880 11008
rect 10692 11024 10744 11076
rect 11980 11024 12032 11076
rect 10416 10956 10468 11008
rect 11336 10956 11388 11008
rect 17132 11024 17184 11076
rect 13452 10956 13504 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 5540 10752 5592 10804
rect 6736 10795 6788 10804
rect 6736 10761 6745 10795
rect 6745 10761 6779 10795
rect 6779 10761 6788 10795
rect 6736 10752 6788 10761
rect 14556 10752 14608 10804
rect 14740 10795 14792 10804
rect 14740 10761 14749 10795
rect 14749 10761 14783 10795
rect 14783 10761 14792 10795
rect 14740 10752 14792 10761
rect 3056 10616 3108 10668
rect 3516 10616 3568 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 7012 10616 7064 10668
rect 10692 10616 10744 10668
rect 12440 10616 12492 10668
rect 13820 10616 13872 10668
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 15108 10616 15160 10668
rect 17592 10616 17644 10668
rect 5724 10548 5776 10600
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 5908 10548 5960 10557
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 14372 10548 14424 10600
rect 14832 10591 14884 10600
rect 14832 10557 14841 10591
rect 14841 10557 14875 10591
rect 14875 10557 14884 10591
rect 14832 10548 14884 10557
rect 4528 10480 4580 10532
rect 848 10412 900 10464
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 8208 10412 8260 10464
rect 10324 10412 10376 10464
rect 11152 10412 11204 10464
rect 12164 10412 12216 10464
rect 12716 10412 12768 10464
rect 16212 10412 16264 10464
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3056 10208 3108 10260
rect 3608 10072 3660 10124
rect 5448 10208 5500 10260
rect 8760 10208 8812 10260
rect 11060 10208 11112 10260
rect 12900 10208 12952 10260
rect 14556 10208 14608 10260
rect 17592 10251 17644 10260
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 5908 10140 5960 10192
rect 6828 10072 6880 10124
rect 9128 10140 9180 10192
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 8484 10072 8536 10124
rect 12716 10140 12768 10192
rect 13268 10140 13320 10192
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 8300 10047 8352 10056
rect 3884 9936 3936 9988
rect 5632 9936 5684 9988
rect 6736 9936 6788 9988
rect 8300 10013 8309 10047
rect 8309 10013 8343 10047
rect 8343 10013 8352 10047
rect 8300 10004 8352 10013
rect 8760 10004 8812 10056
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 5540 9868 5592 9920
rect 6828 9868 6880 9920
rect 11060 10004 11112 10056
rect 11244 10004 11296 10056
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 12164 10004 12216 10056
rect 12624 10004 12676 10056
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 12992 10004 13044 10056
rect 9680 9868 9732 9920
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 12900 9911 12952 9920
rect 12900 9877 12909 9911
rect 12909 9877 12943 9911
rect 12943 9877 12952 9911
rect 12900 9868 12952 9877
rect 13912 10004 13964 10056
rect 15108 10004 15160 10056
rect 15200 10047 15252 10056
rect 15200 10013 15209 10047
rect 15209 10013 15243 10047
rect 15243 10013 15252 10047
rect 15200 10004 15252 10013
rect 15936 10072 15988 10124
rect 16212 10115 16264 10124
rect 16212 10081 16221 10115
rect 16221 10081 16255 10115
rect 16255 10081 16264 10115
rect 16212 10072 16264 10081
rect 13176 9868 13228 9920
rect 16028 9868 16080 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 1768 9664 1820 9716
rect 3884 9707 3936 9716
rect 3884 9673 3893 9707
rect 3893 9673 3927 9707
rect 3927 9673 3936 9707
rect 3884 9664 3936 9673
rect 5632 9664 5684 9716
rect 5816 9707 5868 9716
rect 5816 9673 5825 9707
rect 5825 9673 5859 9707
rect 5859 9673 5868 9707
rect 5816 9664 5868 9673
rect 6736 9664 6788 9716
rect 8484 9664 8536 9716
rect 12716 9664 12768 9716
rect 1676 9596 1728 9648
rect 2136 9571 2188 9580
rect 2136 9537 2151 9571
rect 2151 9537 2185 9571
rect 2185 9537 2188 9571
rect 2136 9528 2188 9537
rect 2964 9528 3016 9580
rect 5540 9528 5592 9580
rect 6828 9596 6880 9648
rect 5908 9528 5960 9580
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3424 9503 3476 9512
rect 3056 9460 3108 9469
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 1584 9392 1636 9444
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 4620 9460 4672 9512
rect 7196 9528 7248 9580
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 8300 9528 8352 9580
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 6552 9460 6604 9512
rect 8484 9460 8536 9512
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 11060 9528 11112 9580
rect 11152 9571 11204 9580
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 11612 9528 11664 9580
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 13268 9707 13320 9716
rect 13268 9673 13277 9707
rect 13277 9673 13311 9707
rect 13311 9673 13320 9707
rect 13268 9664 13320 9673
rect 13360 9707 13412 9716
rect 13360 9673 13369 9707
rect 13369 9673 13403 9707
rect 13403 9673 13412 9707
rect 13360 9664 13412 9673
rect 14556 9707 14608 9716
rect 14556 9673 14565 9707
rect 14565 9673 14599 9707
rect 14599 9673 14608 9707
rect 14556 9664 14608 9673
rect 13912 9528 13964 9580
rect 14924 9639 14976 9648
rect 14924 9605 14933 9639
rect 14933 9605 14967 9639
rect 14967 9605 14976 9639
rect 14924 9596 14976 9605
rect 12716 9460 12768 9469
rect 1952 9324 2004 9376
rect 6920 9392 6972 9444
rect 11796 9392 11848 9444
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 15108 9571 15160 9580
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 13544 9460 13596 9469
rect 17408 9460 17460 9512
rect 6368 9324 6420 9376
rect 11612 9324 11664 9376
rect 12256 9324 12308 9376
rect 12992 9324 13044 9376
rect 14648 9324 14700 9376
rect 17684 9435 17736 9444
rect 17684 9401 17693 9435
rect 17693 9401 17727 9435
rect 17727 9401 17736 9435
rect 17684 9392 17736 9401
rect 14832 9324 14884 9376
rect 15016 9324 15068 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 1584 9120 1636 9172
rect 2964 9120 3016 9172
rect 6368 9163 6420 9172
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 6828 9120 6880 9172
rect 5908 9052 5960 9104
rect 6460 9052 6512 9104
rect 7656 9052 7708 9104
rect 6552 8984 6604 9036
rect 10324 9120 10376 9172
rect 12624 9120 12676 9172
rect 12808 9120 12860 9172
rect 15200 9163 15252 9172
rect 15200 9129 15209 9163
rect 15209 9129 15243 9163
rect 15243 9129 15252 9163
rect 15200 9120 15252 9129
rect 17500 9120 17552 9172
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 14464 9052 14516 9104
rect 10508 8984 10560 9036
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 6828 8916 6880 8968
rect 6460 8848 6512 8900
rect 6736 8848 6788 8900
rect 9220 8916 9272 8968
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 9496 8916 9548 8925
rect 6552 8823 6604 8832
rect 6552 8789 6561 8823
rect 6561 8789 6595 8823
rect 6595 8789 6604 8823
rect 6552 8780 6604 8789
rect 7196 8780 7248 8832
rect 9312 8848 9364 8900
rect 10232 8916 10284 8968
rect 11428 8984 11480 9036
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 15936 9027 15988 9036
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 12256 8916 12308 8968
rect 9772 8891 9824 8900
rect 9772 8857 9781 8891
rect 9781 8857 9815 8891
rect 9815 8857 9824 8891
rect 9772 8848 9824 8857
rect 12900 8916 12952 8968
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 14832 8916 14884 8968
rect 14924 8916 14976 8968
rect 16028 8916 16080 8968
rect 14372 8848 14424 8900
rect 13360 8780 13412 8832
rect 16212 8780 16264 8832
rect 17684 8823 17736 8832
rect 17684 8789 17693 8823
rect 17693 8789 17727 8823
rect 17727 8789 17736 8823
rect 17684 8780 17736 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 7564 8576 7616 8628
rect 8024 8508 8076 8560
rect 9772 8576 9824 8628
rect 11428 8576 11480 8628
rect 10600 8508 10652 8560
rect 1952 8440 2004 8492
rect 3148 8440 3200 8492
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 7932 8440 7984 8492
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 11336 8508 11388 8560
rect 12256 8508 12308 8560
rect 11152 8440 11204 8492
rect 14372 8508 14424 8560
rect 5816 8372 5868 8424
rect 9220 8372 9272 8424
rect 2044 8347 2096 8356
rect 2044 8313 2053 8347
rect 2053 8313 2087 8347
rect 2087 8313 2096 8347
rect 2044 8304 2096 8313
rect 8116 8304 8168 8356
rect 12256 8304 12308 8356
rect 12624 8372 12676 8424
rect 13544 8372 13596 8424
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 17408 8440 17460 8492
rect 15476 8372 15528 8424
rect 16212 8372 16264 8424
rect 14740 8304 14792 8356
rect 14832 8347 14884 8356
rect 14832 8313 14841 8347
rect 14841 8313 14875 8347
rect 14875 8313 14884 8347
rect 14832 8304 14884 8313
rect 17684 8347 17736 8356
rect 17684 8313 17693 8347
rect 17693 8313 17727 8347
rect 17727 8313 17736 8347
rect 17684 8304 17736 8313
rect 1492 8236 1544 8288
rect 3332 8236 3384 8288
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 11980 8279 12032 8288
rect 11980 8245 11989 8279
rect 11989 8245 12023 8279
rect 12023 8245 12032 8279
rect 11980 8236 12032 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3148 8075 3200 8084
rect 3148 8041 3157 8075
rect 3157 8041 3191 8075
rect 3191 8041 3200 8075
rect 3148 8032 3200 8041
rect 5632 8032 5684 8084
rect 7380 8032 7432 8084
rect 9496 8032 9548 8084
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 12992 8075 13044 8084
rect 12992 8041 13001 8075
rect 13001 8041 13035 8075
rect 13035 8041 13044 8075
rect 12992 8032 13044 8041
rect 14832 8032 14884 8084
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 1860 7828 1912 7880
rect 3424 7871 3476 7880
rect 1400 7760 1452 7812
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 6920 7896 6972 7948
rect 3424 7828 3476 7837
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 4804 7828 4856 7880
rect 6552 7871 6604 7880
rect 6552 7837 6570 7871
rect 6570 7837 6604 7871
rect 6552 7828 6604 7837
rect 7748 7828 7800 7880
rect 9404 7964 9456 8016
rect 12532 7964 12584 8016
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 9496 7828 9548 7880
rect 2320 7760 2372 7812
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 10232 7896 10284 7948
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 12072 7896 12124 7948
rect 12992 7896 13044 7948
rect 17408 7939 17460 7948
rect 10968 7760 11020 7812
rect 848 7692 900 7744
rect 3516 7692 3568 7744
rect 8024 7692 8076 7744
rect 10416 7692 10468 7744
rect 14556 7828 14608 7880
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 17408 7905 17417 7939
rect 17417 7905 17451 7939
rect 17451 7905 17460 7939
rect 17408 7896 17460 7905
rect 12532 7692 12584 7744
rect 14188 7692 14240 7744
rect 15752 7692 15804 7744
rect 16764 7735 16816 7744
rect 16764 7701 16773 7735
rect 16773 7701 16807 7735
rect 16807 7701 16816 7735
rect 16764 7692 16816 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1492 7531 1544 7540
rect 1492 7497 1501 7531
rect 1501 7497 1535 7531
rect 1535 7497 1544 7531
rect 1492 7488 1544 7497
rect 2320 7531 2372 7540
rect 2320 7497 2329 7531
rect 2329 7497 2363 7531
rect 2363 7497 2372 7531
rect 2320 7488 2372 7497
rect 4712 7488 4764 7540
rect 5816 7531 5868 7540
rect 5816 7497 5825 7531
rect 5825 7497 5859 7531
rect 5859 7497 5868 7531
rect 5816 7488 5868 7497
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 15752 7531 15804 7540
rect 15752 7497 15761 7531
rect 15761 7497 15795 7531
rect 15795 7497 15804 7531
rect 15752 7488 15804 7497
rect 1860 7420 1912 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 3332 7352 3384 7404
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 6920 7420 6972 7472
rect 7564 7463 7616 7472
rect 7564 7429 7573 7463
rect 7573 7429 7607 7463
rect 7607 7429 7616 7463
rect 7564 7420 7616 7429
rect 10692 7420 10744 7472
rect 4712 7352 4764 7404
rect 5908 7352 5960 7404
rect 7932 7352 7984 7404
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 10416 7352 10468 7404
rect 11336 7352 11388 7404
rect 12072 7420 12124 7472
rect 12256 7463 12308 7472
rect 12256 7429 12265 7463
rect 12265 7429 12299 7463
rect 12299 7429 12308 7463
rect 12256 7420 12308 7429
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 12808 7352 12860 7404
rect 15200 7420 15252 7472
rect 14188 7352 14240 7404
rect 16764 7352 16816 7404
rect 3700 7327 3752 7336
rect 3700 7293 3709 7327
rect 3709 7293 3743 7327
rect 3743 7293 3752 7327
rect 3700 7284 3752 7293
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 10232 7284 10284 7336
rect 5816 7148 5868 7200
rect 7380 7148 7432 7200
rect 7564 7148 7616 7200
rect 11612 7148 11664 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 4712 6944 4764 6996
rect 10324 6944 10376 6996
rect 4160 6876 4212 6928
rect 4620 6876 4672 6928
rect 1584 6808 1636 6860
rect 2780 6808 2832 6860
rect 3608 6808 3660 6860
rect 4068 6808 4120 6860
rect 2136 6740 2188 6792
rect 2964 6740 3016 6792
rect 3332 6740 3384 6792
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 5908 6876 5960 6928
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 10968 6808 11020 6860
rect 11336 6808 11388 6860
rect 1952 6604 2004 6656
rect 3516 6604 3568 6656
rect 6920 6672 6972 6724
rect 8576 6672 8628 6724
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 10416 6740 10468 6792
rect 10600 6783 10652 6792
rect 10600 6749 10609 6783
rect 10609 6749 10643 6783
rect 10643 6749 10652 6783
rect 10600 6740 10652 6749
rect 11612 6740 11664 6792
rect 11980 6808 12032 6860
rect 11888 6740 11940 6792
rect 12072 6740 12124 6792
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 10416 6604 10468 6656
rect 10876 6604 10928 6656
rect 12440 6672 12492 6724
rect 11612 6604 11664 6656
rect 12256 6647 12308 6656
rect 12256 6613 12265 6647
rect 12265 6613 12299 6647
rect 12299 6613 12308 6647
rect 12256 6604 12308 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2136 6400 2188 6452
rect 3516 6400 3568 6452
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 10600 6400 10652 6452
rect 12532 6400 12584 6452
rect 4804 6332 4856 6384
rect 8116 6375 8168 6384
rect 8116 6341 8125 6375
rect 8125 6341 8159 6375
rect 8159 6341 8168 6375
rect 8116 6332 8168 6341
rect 2136 6264 2188 6316
rect 7932 6264 7984 6316
rect 4620 6196 4672 6248
rect 1676 6060 1728 6112
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 3608 6128 3660 6180
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 9956 6332 10008 6384
rect 8392 6196 8444 6248
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 9588 6264 9640 6316
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 3976 6060 4028 6112
rect 4160 6060 4212 6112
rect 6920 6060 6972 6112
rect 9036 6060 9088 6112
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 10508 6060 10560 6112
rect 10784 6060 10836 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 4068 5856 4120 5908
rect 3516 5788 3568 5840
rect 1952 5695 2004 5704
rect 1952 5661 1961 5695
rect 1961 5661 1995 5695
rect 1995 5661 2004 5695
rect 1952 5652 2004 5661
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 3056 5763 3108 5772
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 3056 5720 3108 5729
rect 3700 5720 3752 5772
rect 3976 5720 4028 5772
rect 1676 5584 1728 5636
rect 2780 5652 2832 5704
rect 3516 5652 3568 5704
rect 4804 5856 4856 5908
rect 11980 5856 12032 5908
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 2688 5516 2740 5568
rect 3700 5584 3752 5636
rect 4436 5516 4488 5568
rect 4712 5584 4764 5636
rect 5540 5516 5592 5568
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 6920 5652 6972 5704
rect 7380 5652 7432 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 9312 5652 9364 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 10784 5695 10836 5704
rect 10784 5661 10802 5695
rect 10802 5661 10836 5695
rect 10784 5652 10836 5661
rect 7288 5584 7340 5636
rect 9036 5584 9088 5636
rect 10508 5584 10560 5636
rect 11336 5652 11388 5704
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 11888 5695 11940 5704
rect 11888 5661 11897 5695
rect 11897 5661 11931 5695
rect 11931 5661 11940 5695
rect 11888 5652 11940 5661
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 12348 5652 12400 5704
rect 7104 5516 7156 5568
rect 8300 5516 8352 5568
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 10416 5516 10468 5568
rect 11336 5516 11388 5568
rect 11888 5516 11940 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 3056 5312 3108 5364
rect 4712 5312 4764 5364
rect 6276 5312 6328 5364
rect 8300 5312 8352 5364
rect 2964 5176 3016 5228
rect 3792 5176 3844 5228
rect 7196 5287 7248 5296
rect 7196 5253 7205 5287
rect 7205 5253 7239 5287
rect 7239 5253 7248 5287
rect 7196 5244 7248 5253
rect 7564 5287 7616 5296
rect 7564 5253 7573 5287
rect 7573 5253 7607 5287
rect 7607 5253 7616 5287
rect 7564 5244 7616 5253
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 4436 5176 4488 5228
rect 5816 5176 5868 5228
rect 5908 5176 5960 5228
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 3976 5040 4028 5092
rect 4068 4972 4120 5024
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 4804 5040 4856 5092
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 7104 5040 7156 5092
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 7196 5015 7248 5024
rect 7196 4981 7205 5015
rect 7205 4981 7239 5015
rect 7239 4981 7248 5015
rect 7196 4972 7248 4981
rect 7564 4972 7616 5024
rect 8760 5312 8812 5364
rect 12164 5312 12216 5364
rect 9036 5176 9088 5228
rect 9312 5176 9364 5228
rect 12256 5219 12308 5228
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 12256 5176 12308 5185
rect 12624 5176 12676 5228
rect 8760 5108 8812 5160
rect 9128 5108 9180 5160
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12624 4768 12676 4820
rect 12808 4743 12860 4752
rect 12808 4709 12817 4743
rect 12817 4709 12851 4743
rect 12851 4709 12860 4743
rect 12808 4700 12860 4709
rect 7196 4632 7248 4684
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 10048 4632 10100 4684
rect 12440 4675 12492 4684
rect 12440 4641 12449 4675
rect 12449 4641 12483 4675
rect 12483 4641 12492 4675
rect 12440 4632 12492 4641
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 12256 4564 12308 4616
rect 13636 4564 13688 4616
rect 17776 4607 17828 4616
rect 17776 4573 17785 4607
rect 17785 4573 17819 4607
rect 17819 4573 17828 4607
rect 17776 4564 17828 4573
rect 9956 4496 10008 4548
rect 3976 4428 4028 4480
rect 6092 4428 6144 4480
rect 8760 4471 8812 4480
rect 8760 4437 8769 4471
rect 8769 4437 8803 4471
rect 8803 4437 8812 4471
rect 8760 4428 8812 4437
rect 8944 4471 8996 4480
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 12716 4496 12768 4548
rect 12992 4471 13044 4480
rect 12992 4437 13001 4471
rect 13001 4437 13035 4471
rect 13035 4437 13044 4471
rect 12992 4428 13044 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4620 4224 4672 4276
rect 6644 4224 6696 4276
rect 4068 4156 4120 4208
rect 10048 4267 10100 4276
rect 10048 4233 10057 4267
rect 10057 4233 10091 4267
rect 10091 4233 10100 4267
rect 10048 4224 10100 4233
rect 10784 4224 10836 4276
rect 3976 4088 4028 4140
rect 4804 4088 4856 4140
rect 5908 4088 5960 4140
rect 6092 4131 6144 4140
rect 6092 4097 6101 4131
rect 6101 4097 6135 4131
rect 6135 4097 6144 4131
rect 6092 4088 6144 4097
rect 6736 4131 6788 4140
rect 6736 4097 6745 4131
rect 6745 4097 6779 4131
rect 6779 4097 6788 4131
rect 6736 4088 6788 4097
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 8944 4156 8996 4208
rect 11612 4156 11664 4208
rect 12808 4199 12860 4208
rect 12808 4165 12842 4199
rect 12842 4165 12860 4199
rect 12808 4156 12860 4165
rect 7012 4020 7064 4072
rect 9036 4088 9088 4140
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 7288 3995 7340 4004
rect 7288 3961 7297 3995
rect 7297 3961 7331 3995
rect 7331 3961 7340 3995
rect 7288 3952 7340 3961
rect 4620 3884 4672 3936
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 5356 3884 5408 3936
rect 7012 3884 7064 3936
rect 7104 3884 7156 3936
rect 10508 4020 10560 4072
rect 11060 4063 11112 4072
rect 11060 4029 11069 4063
rect 11069 4029 11103 4063
rect 11103 4029 11112 4063
rect 11060 4020 11112 4029
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 11980 4088 12032 4140
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 11244 3952 11296 4004
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 10232 3884 10284 3936
rect 10508 3884 10560 3936
rect 12256 4020 12308 4072
rect 12440 4020 12492 4072
rect 12348 3884 12400 3936
rect 14004 3927 14056 3936
rect 14004 3893 14013 3927
rect 14013 3893 14047 3927
rect 14047 3893 14056 3927
rect 14004 3884 14056 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 6736 3680 6788 3732
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 10324 3680 10376 3732
rect 12716 3680 12768 3732
rect 12992 3680 13044 3732
rect 4620 3612 4672 3664
rect 5724 3612 5776 3664
rect 9496 3655 9548 3664
rect 9496 3621 9505 3655
rect 9505 3621 9539 3655
rect 9539 3621 9548 3655
rect 9496 3612 9548 3621
rect 9956 3612 10008 3664
rect 11888 3612 11940 3664
rect 12440 3612 12492 3664
rect 7932 3544 7984 3596
rect 4804 3476 4856 3528
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 7380 3476 7432 3528
rect 5816 3408 5868 3460
rect 7840 3476 7892 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 9588 3476 9640 3528
rect 11244 3544 11296 3596
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 11152 3519 11204 3528
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 14004 3476 14056 3528
rect 4528 3383 4580 3392
rect 4528 3349 4537 3383
rect 4537 3349 4571 3383
rect 4571 3349 4580 3383
rect 4528 3340 4580 3349
rect 6460 3340 6512 3392
rect 6920 3340 6972 3392
rect 11060 3408 11112 3460
rect 11612 3408 11664 3460
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 8392 3340 8444 3392
rect 12164 3383 12216 3392
rect 12164 3349 12179 3383
rect 12179 3349 12213 3383
rect 12213 3349 12216 3383
rect 12164 3340 12216 3349
rect 13544 3340 13596 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 6460 3179 6512 3188
rect 6460 3145 6469 3179
rect 6469 3145 6503 3179
rect 6503 3145 6512 3179
rect 6460 3136 6512 3145
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 11060 3136 11112 3188
rect 11612 3179 11664 3188
rect 11612 3145 11621 3179
rect 11621 3145 11655 3179
rect 11655 3145 11664 3179
rect 11612 3136 11664 3145
rect 4528 3068 4580 3120
rect 5724 3000 5776 3052
rect 7196 3068 7248 3120
rect 5540 2932 5592 2984
rect 6828 3000 6880 3052
rect 7840 3068 7892 3120
rect 9496 3111 9548 3120
rect 9496 3077 9530 3111
rect 9530 3077 9548 3111
rect 9496 3068 9548 3077
rect 6920 2932 6972 2984
rect 8576 2975 8628 2984
rect 8576 2941 8585 2975
rect 8585 2941 8619 2975
rect 8619 2941 8628 2975
rect 8576 2932 8628 2941
rect 11152 3111 11204 3120
rect 11152 3077 11161 3111
rect 11161 3077 11195 3111
rect 11195 3077 11204 3111
rect 11152 3068 11204 3077
rect 11244 3000 11296 3052
rect 12624 3136 12676 3188
rect 12532 3068 12584 3120
rect 12164 3000 12216 3052
rect 7380 2864 7432 2916
rect 11888 2932 11940 2984
rect 10784 2907 10836 2916
rect 10784 2873 10793 2907
rect 10793 2873 10827 2907
rect 10827 2873 10836 2907
rect 10784 2864 10836 2873
rect 5908 2796 5960 2848
rect 9404 2796 9456 2848
rect 11152 2796 11204 2848
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 12440 2796 12492 2848
rect 13360 2796 13412 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 13544 2635 13596 2644
rect 13544 2601 13553 2635
rect 13553 2601 13587 2635
rect 13587 2601 13596 2635
rect 13544 2592 13596 2601
rect 8576 2524 8628 2576
rect 7380 2499 7432 2508
rect 7380 2465 7389 2499
rect 7389 2465 7423 2499
rect 7423 2465 7432 2499
rect 7380 2456 7432 2465
rect 5540 2431 5592 2440
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 6828 2388 6880 2440
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 8116 2388 8168 2440
rect 8760 2388 8812 2440
rect 12256 2524 12308 2576
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 11060 2431 11112 2440
rect 11060 2397 11069 2431
rect 11069 2397 11103 2431
rect 11103 2397 11112 2431
rect 11060 2388 11112 2397
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 12072 2388 12124 2440
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 8300 2320 8352 2372
rect 5816 2252 5868 2304
rect 6460 2252 6512 2304
rect 7012 2252 7064 2304
rect 7748 2252 7800 2304
rect 9036 2252 9088 2304
rect 9680 2252 9732 2304
rect 10324 2252 10376 2304
rect 10968 2252 11020 2304
rect 11612 2252 11664 2304
rect 12900 2252 12952 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 8390 20754 8446 21448
rect 9034 20754 9090 21448
rect 10966 20754 11022 21448
rect 8390 20726 8616 20754
rect 8390 20648 8446 20726
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 8588 18970 8616 20726
rect 9034 20726 9260 20754
rect 9034 20648 9090 20726
rect 9232 18970 9260 20726
rect 10888 20726 11022 20754
rect 10888 18970 10916 20726
rect 10966 20648 11022 20726
rect 11610 20754 11666 21448
rect 11610 20726 11928 20754
rect 11610 20648 11666 20726
rect 11900 18970 11928 20726
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 10876 18964 10928 18970
rect 10876 18906 10928 18912
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 848 14544 900 14550
rect 846 14512 848 14521
rect 900 14512 902 14521
rect 846 14447 902 14456
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 4816 14074 4844 14350
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 848 13184 900 13190
rect 846 13152 848 13161
rect 900 13152 902 13161
rect 846 13087 902 13096
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12345 1532 12582
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 848 11552 900 11558
rect 846 11520 848 11529
rect 900 11520 902 11529
rect 846 11455 902 11464
rect 848 10464 900 10470
rect 846 10432 848 10441
rect 900 10432 902 10441
rect 846 10367 902 10376
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1596 9450 1624 9998
rect 1780 9722 1808 9998
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 1688 9330 1716 9590
rect 1596 9302 1716 9330
rect 1596 9178 1624 9302
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1492 8288 1544 8294
rect 1492 8230 1544 8236
rect 1400 7812 1452 7818
rect 1400 7754 1452 7760
rect 848 7744 900 7750
rect 846 7712 848 7721
rect 900 7712 902 7721
rect 846 7647 902 7656
rect 1412 7410 1440 7754
rect 1504 7546 1532 8230
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1596 7342 1624 9114
rect 1872 7886 1900 9998
rect 2148 9586 2176 14010
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12238 4660 13262
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5552 12434 5580 12786
rect 5552 12406 5672 12434
rect 4620 12232 4672 12238
rect 5540 12232 5592 12238
rect 5460 12192 5540 12220
rect 4672 12180 4752 12186
rect 4620 12174 4752 12180
rect 4632 12158 4752 12174
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2976 9586 3004 10406
rect 3068 10266 3096 10610
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1964 8498 1992 9318
rect 2976 9178 3004 9522
rect 3068 9518 3096 10202
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 2056 8265 2084 8298
rect 2042 8256 2098 8265
rect 2042 8191 2098 8200
rect 3160 8090 3188 8434
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 6866 1624 7278
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1688 6118 1716 7822
rect 1872 7478 1900 7822
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2332 7546 2360 7754
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1964 6905 1992 7142
rect 1950 6896 2006 6905
rect 1950 6831 2006 6840
rect 2148 6798 2176 7346
rect 3160 7342 3188 8026
rect 3344 7410 3372 8230
rect 3436 7886 3464 9454
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3528 7834 3556 10610
rect 3620 10130 3648 11630
rect 3896 11354 3924 11698
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 4632 11286 4660 12038
rect 4724 11898 4752 12158
rect 5460 12102 5488 12192
rect 5540 12174 5592 12180
rect 5644 12170 5672 12406
rect 6288 12374 6316 14350
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 13938 6776 14214
rect 8772 14074 8800 18702
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6380 13530 6408 13874
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6380 12442 6408 12854
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6288 12238 6316 12310
rect 6380 12238 6408 12378
rect 6564 12374 6592 13330
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6552 12368 6604 12374
rect 6472 12316 6552 12322
rect 6472 12310 6604 12316
rect 6472 12294 6592 12310
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 5460 11830 5488 12038
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 4724 11150 4752 11290
rect 4528 11144 4580 11150
rect 4528 11086 4580 11092
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4540 10554 4568 11086
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4540 10538 4660 10554
rect 4528 10532 4660 10538
rect 4580 10526 4660 10532
rect 4528 10474 4580 10480
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3896 9722 3924 9930
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 4632 9518 4660 10526
rect 5460 10266 5488 11766
rect 5644 11762 5672 12106
rect 6288 11898 6316 12174
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10810 5580 10950
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5644 9994 5672 11698
rect 5736 11150 5764 11766
rect 6380 11762 6408 12174
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6472 11354 6500 12294
rect 6656 12186 6684 12582
rect 6564 12158 6684 12186
rect 6564 12102 6592 12158
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 5736 10606 5764 11086
rect 6564 10606 6592 11086
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6748 10810 6776 11018
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 5920 10198 5948 10542
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5552 9586 5580 9862
rect 5644 9722 5672 9930
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 3528 7806 3648 7834
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7410 3556 7686
rect 3620 7410 3648 7806
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5642 1716 6054
rect 1964 5710 1992 6598
rect 2148 6458 2176 6734
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2148 5914 2176 6258
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2792 5710 2820 6802
rect 3344 6798 3372 7346
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 2976 5778 3004 6734
rect 3528 6662 3556 7346
rect 3620 6866 3648 7346
rect 3712 7342 3740 9454
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5644 8974 5672 9658
rect 5828 8974 5856 9658
rect 5920 9586 5948 10134
rect 6564 10062 6592 10542
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 6564 9518 6592 9998
rect 6748 9994 6776 10746
rect 6840 10674 6868 10950
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6840 10130 6868 10610
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6748 9722 6776 9930
rect 6840 9926 6868 10066
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 9178 6408 9318
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 6460 9104 6512 9110
rect 6460 9046 6512 9052
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 5644 8090 5672 8910
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4724 7546 4752 7822
rect 4712 7540 4764 7546
rect 4632 7500 4712 7528
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 6458 3556 6598
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 5778 3096 6054
rect 3528 5846 3556 6394
rect 3620 6186 3648 6802
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 2688 5568 2740 5574
rect 2976 5556 3004 5714
rect 2740 5528 3004 5556
rect 2688 5510 2740 5516
rect 2976 5234 3004 5528
rect 3068 5370 3096 5714
rect 3528 5710 3556 5782
rect 3712 5778 3740 7278
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6934 4660 7500
rect 4712 7482 4764 7488
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4724 7002 4752 7346
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5778 4016 6054
rect 4080 5914 4108 6802
rect 4172 6798 4200 6870
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4172 6118 4200 6734
rect 4816 6390 4844 7822
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5828 7546 5856 8366
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5828 7206 5856 7482
rect 5920 7410 5948 9046
rect 6472 8906 6500 9046
rect 6564 9042 6592 9454
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6748 8906 6776 9658
rect 6840 9654 6868 9862
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6840 9178 6868 9590
rect 6932 9450 6960 13806
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7024 12306 7052 13262
rect 7116 12986 7144 13942
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11762 7052 12038
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7024 10674 7052 11698
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7024 10062 7052 10610
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7208 9586 7236 12582
rect 7484 12238 7512 13330
rect 8128 12986 8156 13874
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7484 11354 7512 12174
rect 7668 11898 7696 12718
rect 7760 12646 7788 12718
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 8220 12442 8248 12786
rect 8864 12782 8892 13670
rect 8956 13462 8984 14010
rect 9600 13938 9628 18702
rect 11348 14618 11376 18702
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 9128 13932 9180 13938
rect 9588 13932 9640 13938
rect 9128 13874 9180 13880
rect 9508 13892 9588 13920
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7656 10056 7708 10062
rect 7760 10044 7788 12242
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8206 11792 8262 11801
rect 8206 11727 8208 11736
rect 8260 11727 8262 11736
rect 8208 11698 8260 11704
rect 8312 11626 8340 11834
rect 8404 11830 8432 12174
rect 8956 12170 8984 13398
rect 9140 13326 9168 13874
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9036 12436 9088 12442
rect 9140 12434 9168 13262
rect 9088 12406 9168 12434
rect 9036 12378 9088 12384
rect 8944 12164 8996 12170
rect 8944 12106 8996 12112
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8772 11898 8800 12038
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8680 11626 8708 11766
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7708 10016 7788 10044
rect 7656 9998 7708 10004
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6840 8974 6868 9114
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6564 7886 6592 8774
rect 6932 7954 6960 9386
rect 7668 9110 7696 9998
rect 8220 9586 8248 10406
rect 8772 10266 8800 11834
rect 9048 11762 9076 12378
rect 9232 12102 9260 13262
rect 9324 13190 9352 13738
rect 9508 13326 9536 13892
rect 9588 13874 9640 13880
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 13326 9904 13670
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12986 9444 13126
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9232 11218 9260 11834
rect 9324 11801 9352 12786
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 11830 9444 12038
rect 9508 11898 9536 12922
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9404 11824 9456 11830
rect 9310 11792 9366 11801
rect 9404 11766 9456 11772
rect 9600 11762 9628 12106
rect 9310 11727 9312 11736
rect 9364 11727 9366 11736
rect 9588 11756 9640 11762
rect 9312 11698 9364 11704
rect 9588 11698 9640 11704
rect 9324 11642 9352 11698
rect 9968 11694 9996 13874
rect 10244 13530 10272 14282
rect 11348 14074 11376 14554
rect 11716 14074 11744 18702
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 17682 14376 17738 14385
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9956 11688 10008 11694
rect 9324 11614 9536 11642
rect 9956 11630 10008 11636
rect 10060 11626 10088 11698
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9416 11150 9444 11494
rect 9508 11218 9536 11614
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8312 9586 8340 9998
rect 8496 9722 8524 10066
rect 8772 10062 8800 10202
rect 9140 10198 9168 11086
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 9692 9926 9720 11222
rect 9784 11150 9812 11494
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 9692 9586 9720 9862
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6932 7478 6960 7890
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4632 5710 4660 6190
rect 4816 5914 4844 6326
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3712 5166 3740 5578
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 5234 4476 5510
rect 4724 5370 4752 5578
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3804 5080 3832 5170
rect 3976 5092 4028 5098
rect 3804 5052 3976 5080
rect 3976 5034 4028 5040
rect 3988 4486 4016 5034
rect 4068 5024 4120 5030
rect 4448 5012 4476 5170
rect 5552 5166 5580 5510
rect 5828 5234 5856 7142
rect 5920 6934 5948 7346
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5920 5234 5948 6870
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6932 6118 6960 6666
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6932 5710 6960 6054
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6288 5370 6316 5646
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4448 4984 4660 5012
rect 4068 4966 4120 4972
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3988 4146 4016 4422
rect 4080 4214 4108 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4282 4660 4984
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4816 4146 4844 5034
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3670 4660 3878
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4816 3534 4844 3878
rect 5368 3534 5396 3878
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4540 3126 4568 3334
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 5552 2990 5580 5102
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 4146 6132 4422
rect 6656 4282 6684 5170
rect 7116 5098 7144 5510
rect 7208 5302 7236 8774
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7392 8090 7420 8434
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7206 7420 8026
rect 7576 7478 7604 8570
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 7886 7788 8230
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7944 7546 7972 8434
rect 8036 7750 8064 8502
rect 8128 8362 8156 9522
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8496 9042 8524 9454
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 10244 8974 10272 12718
rect 10336 12646 10364 13874
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10520 12918 10548 13194
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10612 11898 10640 13126
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 9586 10364 10406
rect 10428 10062 10456 10950
rect 10704 10674 10732 11018
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10704 10062 10732 10610
rect 11072 10266 11100 12786
rect 11164 11150 11192 13738
rect 11716 13394 11744 14010
rect 12912 13938 12940 14350
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11532 12306 11560 12854
rect 11716 12850 11744 13126
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11900 12238 11928 13262
rect 12084 12918 12112 13398
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12084 12434 12112 12854
rect 12636 12714 12664 13874
rect 13924 13530 13952 13874
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12084 12406 12204 12434
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11440 12102 11468 12174
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11440 11830 11468 12038
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11624 11762 11652 12038
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11256 11354 11284 11698
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11152 11144 11204 11150
rect 11336 11144 11388 11150
rect 11204 11104 11284 11132
rect 11152 11086 11204 11092
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11164 10146 11192 10406
rect 11072 10118 11192 10146
rect 11256 10146 11284 11104
rect 11336 11086 11388 11092
rect 11348 11014 11376 11086
rect 11992 11082 12020 11698
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11256 10118 11376 10146
rect 11072 10062 11100 10118
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 11060 10056 11112 10062
rect 11244 10056 11296 10062
rect 11060 9998 11112 10004
rect 11164 10016 11244 10044
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10336 9178 10364 9522
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9048 8401 9076 8434
rect 9232 8430 9260 8910
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9220 8424 9272 8430
rect 9034 8392 9090 8401
rect 8116 8356 8168 8362
rect 9220 8366 9272 8372
rect 9034 8327 9090 8336
rect 8116 8298 8168 8304
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7564 7472 7616 7478
rect 7484 7420 7564 7426
rect 7484 7414 7616 7420
rect 7484 7398 7604 7414
rect 7932 7404 7984 7410
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7300 5234 7328 5578
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4690 7236 4966
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7392 4622 7420 5646
rect 7484 5166 7512 7398
rect 8036 7392 8064 7686
rect 7984 7364 8064 7392
rect 7932 7346 7984 7352
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 5302 7604 7142
rect 7944 6322 7972 7346
rect 8128 6390 8156 8298
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8116 6384 8168 6390
rect 8588 6338 8616 6666
rect 8116 6326 8168 6332
rect 8312 6322 8616 6338
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 8312 6316 8628 6322
rect 8312 6310 8576 6316
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7576 5030 7604 5238
rect 7944 5234 7972 6258
rect 8312 5658 8340 6310
rect 8576 6258 8628 6264
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8404 5710 8432 6190
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 8220 5630 8340 5658
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8116 5228 8168 5234
rect 8220 5216 8248 5630
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 5370 8340 5510
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8168 5188 8248 5216
rect 8300 5228 8352 5234
rect 8116 5170 8168 5176
rect 8404 5216 8432 5646
rect 8772 5370 8800 5646
rect 9048 5642 9076 6054
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9048 5234 9076 5578
rect 8352 5188 8432 5216
rect 9036 5228 9088 5234
rect 8300 5170 8352 5176
rect 9036 5170 9088 5176
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 5724 3664 5776 3670
rect 5630 3632 5686 3641
rect 5776 3624 5856 3652
rect 5724 3606 5776 3612
rect 5630 3567 5686 3576
rect 5644 3534 5672 3567
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5736 3058 5764 3470
rect 5828 3466 5856 3624
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5552 2446 5580 2926
rect 5920 2854 5948 4082
rect 6748 3738 6776 4082
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7024 3942 7052 4014
rect 7116 3942 7144 4082
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 7300 3641 7328 3946
rect 7286 3632 7342 3641
rect 7286 3567 7342 3576
rect 7392 3534 7420 4558
rect 7944 3602 7972 5170
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 6472 3194 6500 3334
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5920 2446 5948 2790
rect 6840 2446 6868 2994
rect 6932 2990 6960 3334
rect 7208 3126 7236 3334
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6932 2446 6960 2926
rect 7392 2922 7420 3470
rect 7852 3126 7880 3470
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7392 2514 7420 2858
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 8128 2446 8156 3878
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8312 2378 8340 5170
rect 9140 5166 9168 6258
rect 9232 5556 9260 8366
rect 9324 7886 9352 8842
rect 9508 8090 9536 8910
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9784 8634 9812 8842
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9416 6458 9444 7958
rect 9508 7886 9536 8026
rect 10244 7954 10272 8910
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9404 6452 9456 6458
rect 9324 6412 9404 6440
rect 9324 5710 9352 6412
rect 9404 6394 9456 6400
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9416 5556 9444 5646
rect 9232 5528 9444 5556
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 8772 4486 8800 5102
rect 9324 4622 9352 5170
rect 9416 4622 9444 5528
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8944 4480 8996 4486
rect 9508 4434 9536 7822
rect 9876 7410 9904 7822
rect 9968 7410 9996 7822
rect 10428 7750 10456 9998
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 9042 10548 9522
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10612 8566 10640 9998
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 7410 10456 7686
rect 10612 7528 10640 8502
rect 10520 7500 10640 7528
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9600 6322 9628 6734
rect 9968 6390 9996 7346
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10244 6780 10272 7278
rect 10336 7002 10364 7346
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10428 6798 10456 7346
rect 10324 6792 10376 6798
rect 10244 6752 10324 6780
rect 10324 6734 10376 6740
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 8944 4422 8996 4428
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7012 2304 7064 2310
rect 7748 2304 7800 2310
rect 7064 2264 7144 2292
rect 7012 2246 7064 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 3238 1320 3294 1329
rect 3238 1255 3294 1264
rect 3252 800 3280 1255
rect 5828 800 5856 2246
rect 6472 800 6500 2246
rect 7116 800 7144 2264
rect 7748 2246 7800 2252
rect 7760 800 7788 2246
rect 8404 800 8432 3334
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8588 2582 8616 2926
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8772 2446 8800 4422
rect 8956 4214 8984 4422
rect 9416 4406 9536 4434
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9048 3738 9076 4082
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9140 3194 9168 3470
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9416 2854 9444 4406
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9508 3126 9536 3606
rect 9600 3534 9628 5510
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9968 4146 9996 4490
rect 10060 4282 10088 4626
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9968 3670 9996 4082
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 10244 3534 10272 3878
rect 10336 3738 10364 6734
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6254 10456 6598
rect 10520 6322 10548 7500
rect 10704 7478 10732 9998
rect 11072 9586 11100 9998
rect 11164 9586 11192 10016
rect 11244 9998 11296 10004
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11164 8498 11192 9522
rect 11348 8566 11376 10118
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11624 9586 11652 9998
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11624 9382 11652 9522
rect 11808 9450 11836 9998
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11440 8634 11468 8978
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10980 6866 11008 7754
rect 11348 7410 11376 8502
rect 11440 7954 11468 8570
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11992 7410 12020 8230
rect 12084 7954 12112 11494
rect 12176 11150 12204 12406
rect 12820 12238 12848 12786
rect 13004 12434 13032 13466
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13464 12986 13492 13194
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13004 12406 13124 12434
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12820 11898 12848 12174
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12360 11150 12388 11698
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12176 10470 12204 11086
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12176 9518 12204 9998
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 8974 12296 9318
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12268 8566 12296 8910
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12452 8378 12480 10610
rect 12636 10062 12664 11086
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10198 12756 10406
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12624 10056 12676 10062
rect 12268 8362 12480 8378
rect 12256 8356 12480 8362
rect 12308 8350 12480 8356
rect 12544 10016 12624 10044
rect 12256 8298 12308 8304
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 7478 12112 7890
rect 12268 7478 12296 8298
rect 12544 8022 12572 10016
rect 12624 9998 12676 10004
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12728 9722 12756 9998
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12636 9178 12664 9522
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12728 9042 12756 9454
rect 12820 9178 12848 11698
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12912 9926 12940 10202
rect 13004 10062 13032 12106
rect 13096 11150 13124 12406
rect 13280 12306 13308 12854
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13280 10198 13308 12242
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13268 10192 13320 10198
rect 13320 10152 13400 10180
rect 13268 10134 13320 10140
rect 12992 10056 13044 10062
rect 13044 10016 13308 10044
rect 12992 9998 13044 10004
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13188 9602 13216 9862
rect 13280 9722 13308 10016
rect 13372 9722 13400 10152
rect 13464 10062 13492 10950
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 12912 9586 13216 9602
rect 12900 9580 13216 9586
rect 12952 9574 13216 9580
rect 12900 9522 12952 9528
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12912 8974 12940 9522
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12636 8090 12664 8366
rect 13004 8090 13032 9318
rect 13372 8838 13400 9658
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13556 8430 13584 9454
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12544 7750 12572 7958
rect 13004 7954 13032 8026
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11348 6866 11376 7346
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10612 6458 10640 6734
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10888 6322 10916 6598
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5574 10456 6190
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10520 5642 10548 6054
rect 10796 5710 10824 6054
rect 11348 5710 11376 6802
rect 11624 6798 11652 7142
rect 11992 6866 12020 7346
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12084 6798 12112 7414
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11624 5710 11652 6598
rect 11900 5710 11928 6734
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11888 5704 11940 5710
rect 11992 5658 12020 5850
rect 11940 5652 12020 5658
rect 11888 5646 12020 5652
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 10428 2446 10456 5510
rect 10520 4078 10548 5578
rect 11348 5574 11376 5646
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10520 3942 10548 4014
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10796 2922 10824 4218
rect 11624 4214 11652 5646
rect 11900 5630 12020 5646
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11900 4146 11928 5510
rect 11992 4146 12020 5630
rect 12176 5370 12204 5646
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12268 5234 12296 6598
rect 12348 5704 12400 5710
rect 12452 5658 12480 6666
rect 12544 6458 12572 7686
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12820 6798 12848 7346
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12544 5794 12572 6394
rect 12544 5766 12664 5794
rect 12400 5652 12572 5658
rect 12348 5646 12572 5652
rect 12360 5630 12572 5646
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12268 4622 12296 5170
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12452 4298 12480 4626
rect 12268 4270 12480 4298
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11072 3466 11100 4014
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11256 3602 11284 3946
rect 11900 3670 11928 4082
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11072 3194 11100 3402
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 11072 2446 11100 3130
rect 11164 3126 11192 3470
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11164 2854 11192 3062
rect 11256 3058 11284 3538
rect 11888 3528 11940 3534
rect 11992 3516 12020 4082
rect 12268 4078 12296 4270
rect 12544 4146 12572 5630
rect 12636 5234 12664 5766
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12636 4826 12664 5170
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12360 3534 12388 3878
rect 12452 3670 12480 4014
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 11940 3488 12020 3516
rect 12348 3528 12400 3534
rect 11888 3470 11940 3476
rect 12348 3470 12400 3476
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11624 3194 11652 3402
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11900 2990 11928 3470
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12176 3058 12204 3334
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 11888 2984 11940 2990
rect 11940 2932 12020 2938
rect 11888 2926 12020 2932
rect 11900 2910 12020 2926
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11796 2848 11848 2854
rect 11848 2808 11928 2836
rect 11796 2790 11848 2796
rect 11900 2446 11928 2808
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11888 2440 11940 2446
rect 11992 2428 12020 2910
rect 12452 2854 12480 3606
rect 12544 3126 12572 4082
rect 12636 3534 12664 4762
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12728 3738 12756 4490
rect 12820 4214 12848 4694
rect 13648 4622 13676 13330
rect 14568 13326 14596 14214
rect 16132 14074 16160 14350
rect 17682 14311 17738 14320
rect 17696 14278 17724 14311
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13832 10674 13860 12582
rect 14384 12442 14412 13126
rect 14752 12782 14780 14010
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14936 13530 14964 13874
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14844 12850 14872 13262
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14752 12322 14780 12718
rect 14844 12374 14872 12786
rect 14476 12306 14780 12322
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 15212 12306 15240 13942
rect 14464 12300 14780 12306
rect 14516 12294 14780 12300
rect 14464 12242 14516 12248
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14752 12186 14780 12294
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14832 12232 14884 12238
rect 14752 12180 14832 12186
rect 14752 12174 14884 12180
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 14384 11286 14412 12174
rect 14568 11626 14596 12174
rect 14752 12158 14872 12174
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14568 11354 14596 11562
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14568 11132 14596 11290
rect 14752 11218 14780 12038
rect 14844 11830 14872 12158
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 15304 11762 15332 12174
rect 15488 12170 15516 14010
rect 17696 13705 17724 14010
rect 17682 13696 17738 13705
rect 17682 13631 17738 13640
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14568 11104 14688 11132
rect 14660 11098 14688 11104
rect 14660 11070 14780 11098
rect 14752 10810 14780 11070
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13924 9586 13952 9998
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 14384 8906 14412 10542
rect 14476 9110 14504 10610
rect 14568 10266 14596 10746
rect 14844 10606 14872 11494
rect 14936 11150 14964 11698
rect 15304 11218 15332 11698
rect 15396 11694 15424 12038
rect 15488 11762 15516 12106
rect 15856 11898 15884 13262
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15396 11150 15424 11630
rect 15856 11150 15884 11834
rect 15948 11354 15976 12786
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 16040 12170 16068 12582
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16028 12164 16080 12170
rect 16028 12106 16080 12112
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16132 11286 16160 11698
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 16224 11150 16252 12174
rect 17144 11694 17172 13262
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17328 12345 17356 13126
rect 17512 12782 17540 13262
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17696 13025 17724 13126
rect 17682 13016 17738 13025
rect 17682 12951 17738 12960
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 12442 17540 12718
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17314 12336 17370 12345
rect 17314 12271 17370 12280
rect 17512 12102 17540 12378
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16684 11150 16712 11494
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14568 9722 14596 10202
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 14648 9376 14700 9382
rect 14832 9376 14884 9382
rect 14648 9318 14700 9324
rect 14752 9324 14832 9330
rect 14752 9318 14884 9324
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 14384 8566 14412 8842
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14568 7886 14596 8910
rect 14660 8498 14688 9318
rect 14752 9302 14872 9318
rect 14752 8498 14780 9302
rect 14936 8974 14964 9590
rect 15028 9382 15056 11086
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15120 10062 15148 10610
rect 16224 10470 16252 11086
rect 17144 11082 17172 11630
rect 17788 11354 17816 11630
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 10130 16252 10406
rect 17604 10266 17632 10610
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17696 10305 17724 10406
rect 17682 10296 17738 10305
rect 17592 10260 17644 10266
rect 17682 10231 17738 10240
rect 17592 10202 17644 10208
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15120 9586 15148 9998
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15212 9178 15240 9998
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15948 9042 15976 10066
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 16040 8974 16068 9862
rect 17682 9616 17738 9625
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 17500 9580 17552 9586
rect 17682 9551 17738 9560
rect 17500 9522 17552 9528
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14752 8362 14780 8434
rect 14844 8362 14872 8910
rect 16224 8838 16252 9522
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8430 16252 8774
rect 17420 8498 17448 9454
rect 17512 9178 17540 9522
rect 17696 9450 17724 9551
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17682 8936 17738 8945
rect 17682 8871 17738 8880
rect 17696 8838 17724 8871
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14844 8090 14872 8298
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14200 7410 14228 7686
rect 15212 7478 15240 7822
rect 15488 7546 15516 8366
rect 17420 7954 17448 8434
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17696 8265 17724 8298
rect 17682 8256 17738 8265
rect 17682 8191 17738 8200
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 15764 7546 15792 7686
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 16776 7410 16804 7686
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 13004 3738 13032 4422
rect 17788 4185 17816 4558
rect 17774 4176 17830 4185
rect 17774 4111 17830 4120
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 14016 3534 14044 3878
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 12636 3194 12664 3470
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 12072 2440 12124 2446
rect 11992 2400 12072 2428
rect 11888 2382 11940 2388
rect 12072 2382 12124 2388
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 9048 800 9076 2246
rect 9692 800 9720 2246
rect 10336 800 10364 2246
rect 10980 800 11008 2246
rect 11624 800 11652 2246
rect 12268 800 12296 2518
rect 13372 2446 13400 2790
rect 13556 2650 13584 3334
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12912 800 12940 2246
rect 3238 0 3294 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
<< via2 >>
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 846 14492 848 14512
rect 848 14492 900 14512
rect 900 14492 902 14512
rect 846 14456 902 14492
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 1398 13640 1454 13696
rect 846 13132 848 13152
rect 848 13132 900 13152
rect 900 13132 902 13152
rect 846 13096 902 13132
rect 1490 12280 1546 12336
rect 846 11500 848 11520
rect 848 11500 900 11520
rect 900 11500 902 11520
rect 846 11464 902 11500
rect 846 10412 848 10432
rect 848 10412 900 10432
rect 900 10412 902 10432
rect 846 10376 902 10412
rect 846 7692 848 7712
rect 848 7692 900 7712
rect 900 7692 902 7712
rect 846 7656 902 7692
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 2042 8200 2098 8256
rect 1950 6840 2006 6896
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 8206 11756 8262 11792
rect 8206 11736 8208 11756
rect 8208 11736 8260 11756
rect 8260 11736 8262 11756
rect 9310 11756 9366 11792
rect 9310 11736 9312 11756
rect 9312 11736 9364 11756
rect 9364 11736 9366 11756
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 9034 8336 9090 8392
rect 5630 3576 5686 3632
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 7286 3576 7342 3632
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 3238 1264 3294 1320
rect 17682 14320 17738 14376
rect 17682 13640 17738 13696
rect 17682 12960 17738 13016
rect 17314 12280 17370 12336
rect 17682 10240 17738 10296
rect 17682 9560 17738 9616
rect 17682 8880 17738 8936
rect 17682 8200 17738 8256
rect 17774 4120 17830 4176
<< metal3 >>
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 17677 14378 17743 14381
rect 18504 14378 19304 14408
rect 17677 14376 19304 14378
rect 17677 14320 17682 14376
rect 17738 14320 19304 14376
rect 17677 14318 19304 14320
rect 0 14288 800 14318
rect 17677 14315 17743 14318
rect 18504 14288 19304 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 17677 13698 17743 13701
rect 18504 13698 19304 13728
rect 17677 13696 19304 13698
rect 17677 13640 17682 13696
rect 17738 13640 19304 13696
rect 17677 13638 19304 13640
rect 17677 13635 17743 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 18504 13608 19304 13638
rect 4210 13567 4526 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 17677 13018 17743 13021
rect 18504 13018 19304 13048
rect 17677 13016 19304 13018
rect 17677 12960 17682 13016
rect 17738 12960 19304 13016
rect 17677 12958 19304 12960
rect 0 12928 800 12958
rect 17677 12955 17743 12958
rect 18504 12928 19304 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 17309 12338 17375 12341
rect 18504 12338 19304 12368
rect 17309 12336 19304 12338
rect 17309 12280 17314 12336
rect 17370 12280 19304 12336
rect 17309 12278 19304 12280
rect 17309 12275 17375 12278
rect 18504 12248 19304 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 8201 11794 8267 11797
rect 9305 11794 9371 11797
rect 8201 11792 9371 11794
rect 8201 11736 8206 11792
rect 8262 11736 9310 11792
rect 9366 11736 9371 11792
rect 8201 11734 9371 11736
rect 8201 11731 8267 11734
rect 9305 11731 9371 11734
rect 0 11658 800 11688
rect 0 11568 858 11658
rect 798 11525 858 11568
rect 798 11520 907 11525
rect 798 11464 846 11520
rect 902 11464 907 11520
rect 798 11462 907 11464
rect 841 11459 907 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 17677 10298 17743 10301
rect 18504 10298 19304 10328
rect 17677 10296 19304 10298
rect 17677 10240 17682 10296
rect 17738 10240 19304 10296
rect 17677 10238 19304 10240
rect 0 10208 800 10238
rect 17677 10235 17743 10238
rect 18504 10208 19304 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 17677 9618 17743 9621
rect 18504 9618 19304 9648
rect 17677 9616 19304 9618
rect 17677 9560 17682 9616
rect 17738 9560 19304 9616
rect 17677 9558 19304 9560
rect 17677 9555 17743 9558
rect 18504 9528 19304 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 17677 8938 17743 8941
rect 18504 8938 19304 8968
rect 17677 8936 19304 8938
rect 17677 8880 17682 8936
rect 17738 8880 19304 8936
rect 17677 8878 19304 8880
rect 17677 8875 17743 8878
rect 18504 8848 19304 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 8334 8332 8340 8396
rect 8404 8394 8410 8396
rect 9029 8394 9095 8397
rect 8404 8392 9095 8394
rect 8404 8336 9034 8392
rect 9090 8336 9095 8392
rect 8404 8334 9095 8336
rect 8404 8332 8410 8334
rect 9029 8331 9095 8334
rect 0 8258 800 8288
rect 2037 8258 2103 8261
rect 0 8256 2103 8258
rect 0 8200 2042 8256
rect 2098 8200 2103 8256
rect 0 8198 2103 8200
rect 0 8168 800 8198
rect 2037 8195 2103 8198
rect 17677 8258 17743 8261
rect 18504 8258 19304 8288
rect 17677 8256 19304 8258
rect 17677 8200 17682 8256
rect 17738 8200 19304 8256
rect 17677 8198 19304 8200
rect 17677 8195 17743 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 18504 8168 19304 8198
rect 4210 8127 4526 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 0 7488 800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 1945 6898 2011 6901
rect 0 6896 2011 6898
rect 0 6840 1950 6896
rect 2006 6840 2011 6896
rect 0 6838 2011 6840
rect 0 6808 800 6838
rect 1945 6835 2011 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 17769 4178 17835 4181
rect 18504 4178 19304 4208
rect 17769 4176 19304 4178
rect 17769 4120 17774 4176
rect 17830 4120 19304 4176
rect 17769 4118 19304 4120
rect 17769 4115 17835 4118
rect 18504 4088 19304 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 5625 3634 5691 3637
rect 7281 3634 7347 3637
rect 5625 3632 7347 3634
rect 5625 3576 5630 3632
rect 5686 3576 7286 3632
rect 7342 3576 7347 3632
rect 5625 3574 7347 3576
rect 5625 3571 5691 3574
rect 7281 3571 7347 3574
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 3233 1322 3299 1325
rect 8334 1322 8340 1324
rect 3233 1320 8340 1322
rect 3233 1264 3238 1320
rect 3294 1264 8340 1320
rect 3233 1262 8340 1264
rect 3233 1259 3299 1262
rect 8334 1260 8340 1262
rect 8404 1260 8410 1324
<< via3 >>
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 8340 8332 8404 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 8340 1260 8404 1324
<< metal4 >>
rect 4208 19072 4528 19088
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 18528 5188 19088
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 8339 8396 8405 8397
rect 8339 8332 8340 8396
rect 8404 8332 8405 8396
rect 8339 8331 8405 8332
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 8342 1325 8402 8331
rect 8339 1324 8405 1325
rect 8339 1260 8340 1324
rect 8404 1260 8405 1324
rect 8339 1259 8405 1260
use sky130_fd_sc_hd__nand2_1  _168_
timestamp 0
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  _169_
timestamp 0
transform 1 0 8280 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _170_
timestamp 0
transform 1 0 9752 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _171_
timestamp 0
transform 1 0 9292 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _172_
timestamp 0
transform -1 0 15088 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _173_
timestamp 0
transform 1 0 15088 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _174_
timestamp 0
transform -1 0 16192 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _175_
timestamp 0
transform -1 0 14996 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _176_
timestamp 0
transform 1 0 14168 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_4  _177_
timestamp 0
transform -1 0 16560 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _178_
timestamp 0
transform -1 0 11776 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _179_
timestamp 0
transform 1 0 11592 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _180_
timestamp 0
transform 1 0 5152 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _181_
timestamp 0
transform 1 0 6256 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_2  _182_
timestamp 0
transform 1 0 5336 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _183_
timestamp 0
transform -1 0 9016 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _184_
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _185_
timestamp 0
transform -1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _186_
timestamp 0
transform -1 0 10028 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _187_
timestamp 0
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_2  _188_
timestamp 0
transform -1 0 9936 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _189_
timestamp 0
transform 1 0 9016 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _190_
timestamp 0
transform 1 0 9568 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _191_
timestamp 0
transform 1 0 9568 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _192_
timestamp 0
transform -1 0 10028 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _193_
timestamp 0
transform -1 0 11316 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _194_
timestamp 0
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _195_
timestamp 0
transform -1 0 11868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _196_
timestamp 0
transform 1 0 9108 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _197_
timestamp 0
transform -1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_2  _198_
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _199_
timestamp 0
transform 1 0 3220 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _200_
timestamp 0
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _201_
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _202_
timestamp 0
transform 1 0 3220 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _203_
timestamp 0
transform -1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _204_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _205_
timestamp 0
transform 1 0 2300 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _206_
timestamp 0
transform -1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 0
transform -1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _208_
timestamp 0
transform 1 0 2760 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _209_
timestamp 0
transform -1 0 2208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _210_
timestamp 0
transform 1 0 3496 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _211_
timestamp 0
transform -1 0 4600 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _212_
timestamp 0
transform 1 0 4324 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _213_
timestamp 0
transform -1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _214_
timestamp 0
transform 1 0 4140 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _215_
timestamp 0
transform -1 0 6164 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _216_
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _217_
timestamp 0
transform -1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _218_
timestamp 0
transform -1 0 6808 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _219_
timestamp 0
transform -1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _220_
timestamp 0
transform -1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _221_
timestamp 0
transform 1 0 9476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _222_
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _223_
timestamp 0
transform -1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _224_
timestamp 0
transform 1 0 11500 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _225_
timestamp 0
transform 1 0 11500 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _226_
timestamp 0
transform 1 0 12052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _227_
timestamp 0
transform -1 0 12512 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _228_
timestamp 0
transform -1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _229_
timestamp 0
transform -1 0 11960 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _230_
timestamp 0
transform -1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _231_
timestamp 0
transform 1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _232_
timestamp 0
transform 1 0 9936 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _233_
timestamp 0
transform -1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _234_
timestamp 0
transform 1 0 12052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _235_
timestamp 0
transform 1 0 11040 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _236_
timestamp 0
transform -1 0 9660 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _237_
timestamp 0
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _238_
timestamp 0
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _239_
timestamp 0
transform 1 0 7544 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _240_
timestamp 0
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _241_
timestamp 0
transform 1 0 9292 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _242_
timestamp 0
transform 1 0 10120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _243_
timestamp 0
transform 1 0 10304 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _244_
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _245_
timestamp 0
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _246_
timestamp 0
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _247_
timestamp 0
transform -1 0 7728 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _248_
timestamp 0
transform 1 0 8188 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _249_
timestamp 0
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _250_
timestamp 0
transform -1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _251_
timestamp 0
transform -1 0 11592 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _252_
timestamp 0
transform -1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _253_
timestamp 0
transform 1 0 8096 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _254_
timestamp 0
transform -1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _255_
timestamp 0
transform -1 0 6164 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _256_
timestamp 0
transform 1 0 5612 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _257_
timestamp 0
transform 1 0 6164 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a41oi_1  _258_
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _259_
timestamp 0
transform 1 0 5520 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _260_
timestamp 0
transform -1 0 5796 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_1  _261_
timestamp 0
transform 1 0 3864 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 0
transform -1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _263_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _264_
timestamp 0
transform 1 0 6808 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _265_
timestamp 0
transform 1 0 4140 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _266_
timestamp 0
transform 1 0 6992 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _267_
timestamp 0
transform -1 0 6992 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _268_
timestamp 0
transform -1 0 7084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _269_
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _270_
timestamp 0
transform 1 0 8188 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _271_
timestamp 0
transform -1 0 8188 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a41oi_1  _272_
timestamp 0
transform -1 0 8004 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _273_
timestamp 0
transform -1 0 7636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _274_
timestamp 0
transform 1 0 8004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _275_
timestamp 0
transform -1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _276_
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _277_
timestamp 0
transform 1 0 9292 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _278_
timestamp 0
transform -1 0 10580 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_2  _279_
timestamp 0
transform 1 0 10304 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _280_
timestamp 0
transform -1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _281_
timestamp 0
transform -1 0 13156 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _282_
timestamp 0
transform -1 0 11132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _283_
timestamp 0
transform -1 0 12696 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _284_
timestamp 0
transform 1 0 13156 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _285_
timestamp 0
transform 1 0 12788 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_2  _286_
timestamp 0
transform 1 0 14076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _287_
timestamp 0
transform -1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _288_
timestamp 0
transform -1 0 14812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _289_
timestamp 0
transform -1 0 15272 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _290_
timestamp 0
transform 1 0 12696 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _291_
timestamp 0
transform -1 0 12512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _292_
timestamp 0
transform 1 0 14996 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _293_
timestamp 0
transform 1 0 14536 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _294_
timestamp 0
transform 1 0 12512 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_1  _295_
timestamp 0
transform -1 0 12972 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _296_
timestamp 0
transform 1 0 14444 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _297_
timestamp 0
transform 1 0 12052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _298_
timestamp 0
transform -1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _299_
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _300_
timestamp 0
transform 1 0 12788 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _301_
timestamp 0
transform 1 0 13432 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _302_
timestamp 0
transform 1 0 12880 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 0
transform -1 0 15088 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _304_
timestamp 0
transform -1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _305_
timestamp 0
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _306_
timestamp 0
transform 1 0 15364 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _307_
timestamp 0
transform -1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _308_
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 0
transform -1 0 16376 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 0
transform -1 0 14996 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 0
transform -1 0 13892 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 0
transform -1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 0
transform -1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 0
transform -1 0 8464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 0
transform 1 0 6716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 0
transform -1 0 4600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 0
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 0
transform -1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 0
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 0
transform -1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 0
transform -1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 0
transform -1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 0
transform 1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 0
transform 1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _326_
timestamp 0
transform -1 0 3680 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _327_
timestamp 0
transform -1 0 3496 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_4  _328_
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _329_
timestamp 0
transform -1 0 8372 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_4  _330_
timestamp 0
transform 1 0 6716 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_4  _331_
timestamp 0
transform -1 0 11040 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _332_
timestamp 0
transform -1 0 12420 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _333_
timestamp 0
transform -1 0 11224 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_4  _334_
timestamp 0
transform -1 0 12052 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _335_
timestamp 0
transform -1 0 8188 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _336_
timestamp 0
transform 1 0 1840 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _337_
timestamp 0
transform 1 0 1748 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _338_
timestamp 0
transform 1 0 4140 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _339_
timestamp 0
transform -1 0 3036 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _340_
timestamp 0
transform 1 0 4600 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _341_
timestamp 0
transform 1 0 3864 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _342_
timestamp 0
transform 1 0 5704 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _343_
timestamp 0
transform 1 0 7360 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _344_
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _345_
timestamp 0
transform 1 0 12512 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _346_
timestamp 0
transform -1 0 13248 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _347_
timestamp 0
transform 1 0 9200 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _348_
timestamp 0
transform 1 0 7176 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _349_
timestamp 0
transform -1 0 11132 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _350_
timestamp 0
transform 1 0 6348 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _351_
timestamp 0
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _352_
timestamp 0
transform -1 0 6900 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _353_
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _354_
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _355_
timestamp 0
transform -1 0 6256 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _356_
timestamp 0
transform -1 0 10396 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _357_
timestamp 0
transform 1 0 7360 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _358_
timestamp 0
transform 1 0 9936 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _359_
timestamp 0
transform -1 0 12972 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _360_
timestamp 0
transform 1 0 14076 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _361_
timestamp 0
transform 1 0 15180 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _362_
timestamp 0
transform 1 0 15916 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _363_
timestamp 0
transform 1 0 16192 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _364_
timestamp 0
transform 1 0 13340 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _365_
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _366_
timestamp 0
transform 1 0 16192 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _367_
timestamp 0
transform 1 0 16376 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 9016 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 8188 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform -1 0 8188 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform 1 0 12236 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 0
transform -1 0 6808 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload1
timestamp 0
transform 1 0 12604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 0
transform -1 0 3220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 0
transform 1 0 10488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 0
transform -1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 0
transform -1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 0
transform 1 0 13156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout44
timestamp 0
transform -1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 0
transform -1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 0
transform -1 0 10396 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 0
transform 1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47
timestamp 0
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91
timestamp 0
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98
timestamp 0
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_105
timestamp 0
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 0
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 0
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 0
transform 1 0 6624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78
timestamp 0
transform 1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_104
timestamp 0
transform 1 0 10672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 0
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_132
timestamp 0
transform 1 0 13248 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_144
timestamp 0
transform 1 0 14352 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_156
timestamp 0
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_35
timestamp 0
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_39
timestamp 0
transform 1 0 4692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_45
timestamp 0
transform 1 0 5244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_79
timestamp 0
transform 1 0 8372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_88
timestamp 0
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_95
timestamp 0
transform 1 0 9844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_100
timestamp 0
transform 1 0 10304 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 0
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 0
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_181
timestamp 0
transform 1 0 17756 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_38
timestamp 0
transform 1 0 4600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_77
timestamp 0
transform 1 0 8188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_89
timestamp 0
transform 1 0 9292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_95
timestamp 0
transform 1 0 9844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 0
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 0
transform 1 0 12420 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_148
timestamp 0
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 0
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_92
timestamp 0
transform 1 0 9568 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_104
timestamp 0
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_116
timestamp 0
transform 1 0 11776 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_122
timestamp 0
transform 1 0 12328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 0
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 0
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_177
timestamp 0
transform 1 0 17388 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_23
timestamp 0
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 0
transform 1 0 3956 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 0
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_90
timestamp 0
transform 1 0 9384 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_102
timestamp 0
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 0
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_124
timestamp 0
transform 1 0 12512 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_136
timestamp 0
transform 1 0 13616 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_148
timestamp 0
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 0
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_181
timestamp 0
transform 1 0 17756 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 0
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_12
timestamp 0
transform 1 0 2208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 0
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 0
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 0
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_177
timestamp 0
transform 1 0 17388 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_181
timestamp 0
transform 1 0 17756 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_26
timestamp 0
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_38
timestamp 0
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 0
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_77
timestamp 0
transform 1 0 8188 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_88
timestamp 0
transform 1 0 9200 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 0
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 0
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_18
timestamp 0
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 0
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_34
timestamp 0
transform 1 0 4232 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_62
timestamp 0
transform 1 0 6808 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_74
timestamp 0
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 0
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 0
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_95
timestamp 0
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_101
timestamp 0
transform 1 0 10396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_106
timestamp 0
transform 1 0 10856 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_112
timestamp 0
transform 1 0 11408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 0
transform 1 0 11868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 0
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 0
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp 0
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp 0
transform 1 0 17756 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_30
timestamp 0
transform 1 0 3864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_49
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 0
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_75
timestamp 0
transform 1 0 8004 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_87
timestamp 0
transform 1 0 9108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 0
transform 1 0 10212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_104
timestamp 0
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 0
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 0
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_63
timestamp 0
transform 1 0 6900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 0
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_113
timestamp 0
transform 1 0 11500 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_119
timestamp 0
transform 1 0 12052 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_126
timestamp 0
transform 1 0 12696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_132
timestamp 0
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 0
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_13
timestamp 0
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_25
timestamp 0
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_37
timestamp 0
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 0
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_65
timestamp 0
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_76
timestamp 0
transform 1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 0
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 0
transform 1 0 10856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_119
timestamp 0
transform 1 0 12052 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_131
timestamp 0
transform 1 0 13156 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 0
transform 1 0 13892 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_153
timestamp 0
transform 1 0 15180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 0
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_177
timestamp 0
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 0
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_60
timestamp 0
transform 1 0 6624 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_72
timestamp 0
transform 1 0 7728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_95
timestamp 0
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp 0
transform 1 0 10212 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_108
timestamp 0
transform 1 0 11040 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 0
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_129
timestamp 0
transform 1 0 12972 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 0
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 0
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_154
timestamp 0
transform 1 0 15272 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_160
timestamp 0
transform 1 0 15824 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_177
timestamp 0
transform 1 0 17388 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_36
timestamp 0
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_48
timestamp 0
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 0
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_80
timestamp 0
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_97
timestamp 0
transform 1 0 10028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 0
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_136
timestamp 0
transform 1 0 13616 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_177
timestamp 0
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 0
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_60
timestamp 0
transform 1 0 6624 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 0
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_119
timestamp 0
transform 1 0 12052 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_125
timestamp 0
transform 1 0 12604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 0
transform 1 0 13524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 0
transform 1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 0
transform 1 0 15272 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_162
timestamp 0
transform 1 0 16008 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_180
timestamp 0
transform 1 0 17664 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_7
timestamp 0
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 0
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 0
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_47
timestamp 0
transform 1 0 5428 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 0
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_64
timestamp 0
transform 1 0 6992 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_76
timestamp 0
transform 1 0 8096 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_88
timestamp 0
transform 1 0 9200 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_100
timestamp 0
transform 1 0 10304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 0
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_150
timestamp 0
transform 1 0 14904 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 0
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_177
timestamp 0
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_44
timestamp 0
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 0
transform 1 0 5796 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_59
timestamp 0
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_66
timestamp 0
transform 1 0 7176 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_78
timestamp 0
transform 1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_100
timestamp 0
transform 1 0 10304 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_108
timestamp 0
transform 1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_114
timestamp 0
transform 1 0 11592 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_118
timestamp 0
transform 1 0 11960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_123
timestamp 0
transform 1 0 12420 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 0
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 0
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 0
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_153
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_161
timestamp 0
transform 1 0 15916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_7
timestamp 0
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_19
timestamp 0
transform 1 0 2852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 0
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 0
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_64
timestamp 0
transform 1 0 6992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp 0
transform 1 0 8096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_86
timestamp 0
transform 1 0 9016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_97
timestamp 0
transform 1 0 10028 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 0
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 0
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_130
timestamp 0
transform 1 0 13064 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 0
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_146
timestamp 0
transform 1 0 14536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_175
timestamp 0
transform 1 0 17204 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 0
transform 1 0 17756 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_38
timestamp 0
transform 1 0 4600 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_64
timestamp 0
transform 1 0 6992 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_71
timestamp 0
transform 1 0 7636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_91
timestamp 0
transform 1 0 9476 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_103
timestamp 0
transform 1 0 10580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_120
timestamp 0
transform 1 0 12144 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_155
timestamp 0
transform 1 0 15364 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 0
transform 1 0 16100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 0
transform 1 0 17664 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_7
timestamp 0
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_19
timestamp 0
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_31
timestamp 0
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_43
timestamp 0
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_67
timestamp 0
transform 1 0 7268 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_78
timestamp 0
transform 1 0 8280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_86
timestamp 0
transform 1 0 9016 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_94
timestamp 0
transform 1 0 9752 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_102
timestamp 0
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 0
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_116
timestamp 0
transform 1 0 11776 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_124
timestamp 0
transform 1 0 12512 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_132
timestamp 0
transform 1 0 13248 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_144
timestamp 0
transform 1 0 14352 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_156
timestamp 0
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 0
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_180
timestamp 0
transform 1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_7
timestamp 0
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 0
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 0
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 0
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_103
timestamp 0
transform 1 0 10580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_111
timestamp 0
transform 1 0 11316 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_122
timestamp 0
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_152
timestamp 0
transform 1 0 15088 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_164
timestamp 0
transform 1 0 16192 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_172
timestamp 0
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_6
timestamp 0
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_18
timestamp 0
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_30
timestamp 0
transform 1 0 3864 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_38
timestamp 0
transform 1 0 4600 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_64
timestamp 0
transform 1 0 6992 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_101
timestamp 0
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 0
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_129
timestamp 0
transform 1 0 12972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 0
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_177
timestamp 0
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_7
timestamp 0
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 0
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_49
timestamp 0
transform 1 0 5612 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_59
timestamp 0
transform 1 0 6532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_71
timestamp 0
transform 1 0 7636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 0
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_112
timestamp 0
transform 1 0 11408 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_124
timestamp 0
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 0
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 0
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_151
timestamp 0
transform 1 0 14996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 0
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_177
timestamp 0
transform 1 0 17388 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 0
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 0
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 0
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_177
timestamp 0
transform 1 0 17388 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_181
timestamp 0
transform 1 0 17756 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 0
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 0
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 0
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 0
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 0
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 0
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 0
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 0
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 0
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_177
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_181
timestamp 0
transform 1 0 17756 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 0
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 0
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 0
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 0
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 0
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 0
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 0
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 0
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 0
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 0
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 0
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 0
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 0
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 0
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 0
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_177
timestamp 0
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_181
timestamp 0
transform 1 0 17756 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 0
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 0
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 0
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 0
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 0
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 0
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 0
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 0
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_181
timestamp 0
transform 1 0 17756 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 0
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 0
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_53
timestamp 0
transform 1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_57
timestamp 0
transform 1 0 6348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_69
timestamp 0
transform 1 0 7452 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_77
timestamp 0
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_91
timestamp 0
transform 1 0 9476 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_103
timestamp 0
transform 1 0 10580 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_107
timestamp 0
transform 1 0 10948 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_113
timestamp 0
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_119
timestamp 0
transform 1 0 12052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 0
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 0
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_165
timestamp 0
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_169
timestamp 0
transform 1 0 16652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_181
timestamp 0
transform 1 0 17756 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 9384 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 11132 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform 1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform -1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform 1 0 5796 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform -1 0 16284 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform -1 0 8556 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform -1 0 14720 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 3220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform -1 0 9568 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform -1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform -1 0 17664 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform -1 0 3220 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 5704 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform 1 0 11592 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform -1 0 5704 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 0
transform 1 0 5244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform 1 0 17572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap38
timestamp 0
transform -1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  max_cap39
timestamp 0
transform 1 0 10672 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap40
timestamp 0
transform 1 0 10304 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 0
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 0
transform -1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 0
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 0
transform -1 0 8832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 0
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 0
transform -1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform -1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform -1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform -1 0 8832 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 0
transform -1 0 11408 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 0
transform 1 0 11684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 0
transform 1 0 17480 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 0
transform 1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 0
transform 1 0 17480 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 0
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 0
transform 1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 0
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 0
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 0
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 0
transform 1 0 17112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 0
transform -1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 0
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 0
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 0
transform -1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 0
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 0
transform -1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 0
transform -1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_31
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_32
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_33
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_34
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_35
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_36
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_37
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_38
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_39
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 18124 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_40
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_41
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_42
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 18124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_43
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_44
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_45
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_46
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_47
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_48
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 18124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_49
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 18124 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_50
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 18124 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_51
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 18124 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_52
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_53
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_54
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 18124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_55
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_56
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 18124 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_57
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 18124 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_58
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 18124 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_59
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 18124 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_60
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 18124 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_61
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 18124 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_68
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_69
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_70
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_71
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_72
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_73
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_74
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_75
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_76
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_78
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_79
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_81
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_82
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_87
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_92
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_93
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_96
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_97
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_101
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_102
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_103
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_104
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_105
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_106
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_107
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_108
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_109
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_110
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_111
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_112
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_113
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_114
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_115
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_116
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_117
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_118
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_119
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_120
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_121
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_122
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_123
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_124
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_125
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_126
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_127
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_128
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_129
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_130
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_131
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_132
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_133
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_134
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_135
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_136
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_137
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_138
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_139
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_140
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_141
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_142
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_143
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_144
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_145
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_146
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_147
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_148
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_151
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_152
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_153
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_154
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_155
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_156
timestamp 0
transform 1 0 6256 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_157
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_158
timestamp 0
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_159
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_160
timestamp 0
transform 1 0 16560 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire37
timestamp 0
transform -1 0 13064 0 -1 11968
box -38 -48 314 592
<< labels >>
rlabel metal1 s 9614 18496 9614 18496 4 VGND
rlabel metal1 s 9614 19040 9614 19040 4 VPWR
rlabel metal1 s 1916 9962 1916 9962 4 _000_
rlabel metal2 s 2346 7650 2346 7650 4 _001_
rlabel metal1 s 4646 6970 4646 6970 4 _002_
rlabel metal1 s 2442 6290 2442 6290 4 _003_
rlabel metal1 s 4462 5338 4462 5338 4 _004_
rlabel metal1 s 4365 3094 4365 3094 4 _005_
rlabel metal1 s 5918 3434 5918 3434 4 _006_
rlabel metal1 s 7907 2414 7907 2414 4 _007_
rlabel metal1 s 12473 5610 12473 5610 4 _008_
rlabel metal2 s 12829 4182 12829 4182 4 _009_
rlabel metal2 s 12190 3196 12190 3196 4 _010_
rlabel metal2 s 9517 3094 9517 3094 4 _011_
rlabel metal1 s 7631 7854 7631 7854 4 _012_
rlabel metal2 s 10814 5678 10814 5678 4 _013_
rlabel metal1 s 6424 5610 6424 5610 4 _014_
rlabel metal1 s 7580 4590 7580 4590 4 _015_
rlabel metal2 s 6582 7854 6582 7854 4 _016_
rlabel metal2 s 3910 9826 3910 9826 4 _017_
rlabel metal1 s 4048 11322 4048 11322 4 _018_
rlabel metal1 s 6087 13974 6087 13974 4 _019_
rlabel metal1 s 9112 9962 9112 9962 4 _020_
rlabel metal2 s 8142 13430 8142 13430 4 _021_
rlabel metal1 s 10212 13498 10212 13498 4 _022_
rlabel metal1 s 11868 12682 11868 12682 4 _023_
rlabel metal1 s 14296 7378 14296 7378 4 _024_
rlabel metal1 s 15400 7854 15400 7854 4 _025_
rlabel metal1 s 16136 8942 16136 8942 4 _026_
rlabel metal1 s 15906 10030 15906 10030 4 _027_
rlabel metal1 s 13892 13498 13892 13498 4 _028_
rlabel metal1 s 15032 13906 15032 13906 4 _029_
rlabel metal1 s 16268 12138 16268 12138 4 _030_
rlabel metal2 s 16693 11118 16693 11118 4 _031_
rlabel metal2 s 14858 11050 14858 11050 4 _032_
rlabel metal2 s 14582 10234 14582 10234 4 _033_
rlabel metal1 s 12834 9486 12834 9486 4 _034_
rlabel metal2 s 14766 8398 14766 8398 4 _035_
rlabel metal1 s 9062 11152 9062 11152 4 _036_
rlabel metal1 s 12558 6800 12558 6800 4 _037_
rlabel metal1 s 6164 11798 6164 11798 4 _038_
rlabel metal1 s 10166 11118 10166 11118 4 _039_
rlabel metal1 s 9614 13260 9614 13260 4 _040_
rlabel metal1 s 9706 11084 9706 11084 4 _041_
rlabel metal1 s 7314 11866 7314 11866 4 _042_
rlabel metal1 s 10350 11764 10350 11764 4 _043_
rlabel metal2 s 9798 11322 9798 11322 4 _044_
rlabel metal1 s 12558 11152 12558 11152 4 _045_
rlabel metal1 s 7406 10132 7406 10132 4 _046_
rlabel metal2 s 11454 12002 11454 12002 4 _047_
rlabel metal2 s 9890 13498 9890 13498 4 _048_
rlabel metal1 s 12512 12886 12512 12886 4 _049_
rlabel metal2 s 8510 9248 8510 9248 4 _050_
rlabel metal2 s 10534 6902 10534 6902 4 _051_
rlabel metal2 s 11638 11900 11638 11900 4 _052_
rlabel metal1 s 12926 10030 12926 10030 4 _053_
rlabel metal1 s 8556 12886 8556 12886 4 _054_
rlabel metal1 s 1840 9418 1840 9418 4 _055_
rlabel metal1 s 14858 7854 14858 7854 4 _056_
rlabel metal2 s 1794 9860 1794 9860 4 _057_
rlabel metal1 s 2254 7344 2254 7344 4 _058_
rlabel metal1 s 3266 7344 3266 7344 4 _059_
rlabel metal1 s 4370 6732 4370 6732 4 _060_
rlabel metal1 s 1886 5746 1886 5746 4 _061_
rlabel metal1 s 4554 6732 4554 6732 4 _062_
rlabel metal1 s 2806 5576 2806 5576 4 _063_
rlabel metal1 s 4094 5168 4094 5168 4 _064_
rlabel metal1 s 4554 5202 4554 5202 4 _065_
rlabel metal1 s 4324 5202 4324 5202 4 _066_
rlabel metal1 s 4462 3536 4462 3536 4 _067_
rlabel metal2 s 5382 3706 5382 3706 4 _068_
rlabel metal1 s 4738 3502 4738 3502 4 _069_
rlabel metal1 s 7222 4080 7222 4080 4 _070_
rlabel metal2 s 5658 3553 5658 3553 4 _071_
rlabel metal1 s 10718 8976 10718 8976 4 _072_
rlabel metal1 s 8556 4182 8556 4182 4 _073_
rlabel metal1 s 12006 5712 12006 5712 4 _074_
rlabel metal1 s 11960 6902 11960 6902 4 _075_
rlabel metal2 s 12282 5916 12282 5916 4 _076_
rlabel metal1 s 12236 5338 12236 5338 4 _077_
rlabel metal2 s 12374 3706 12374 3706 4 _078_
rlabel metal1 s 12788 4522 12788 4522 4 _079_
rlabel metal1 s 10672 3978 10672 3978 4 _080_
rlabel metal2 s 11638 3298 11638 3298 4 _081_
rlabel metal1 s 9246 7922 9246 7922 4 _082_
rlabel metal1 s 9568 3502 9568 3502 4 _083_
rlabel metal1 s 7774 8330 7774 8330 4 _084_
rlabel metal2 s 7958 7990 7958 7990 4 _085_
rlabel metal1 s 11086 6222 11086 6222 4 _086_
rlabel metal1 s 10258 6970 10258 6970 4 _087_
rlabel metal1 s 11086 7174 11086 7174 4 _088_
rlabel metal1 s 11224 6766 11224 6766 4 _089_
rlabel metal2 s 10902 6460 10902 6460 4 _090_
rlabel metal1 s 7222 5066 7222 5066 4 _091_
rlabel metal1 s 6946 5168 6946 5168 4 _092_
rlabel metal1 s 6532 5338 6532 5338 4 _093_
rlabel metal2 s 11270 11526 11270 11526 4 _094_
rlabel metal1 s 7222 13362 7222 13362 4 _095_
rlabel metal2 s 7222 7038 7222 7038 4 _096_
rlabel metal1 s 6210 8840 6210 8840 4 _097_
rlabel metal2 s 6394 9248 6394 9248 4 _098_
rlabel metal1 s 5796 9894 5796 9894 4 _099_
rlabel metal2 s 4554 10812 4554 10812 4 _100_
rlabel metal1 s 5106 11152 5106 11152 4 _101_
rlabel metal1 s 4830 11084 4830 11084 4 _102_
rlabel metal1 s 6808 12818 6808 12818 4 _103_
rlabel metal1 s 6670 13940 6670 13940 4 _104_
rlabel metal1 s 7774 9996 7774 9996 4 _105_
rlabel metal2 s 8234 9996 8234 9996 4 _106_
rlabel metal1 s 6624 13498 6624 13498 4 _107_
rlabel metal1 s 8464 9690 8464 9690 4 _108_
rlabel metal1 s 8004 12818 8004 12818 4 _109_
rlabel metal1 s 7820 12410 7820 12410 4 _110_
rlabel metal1 s 10480 13158 10480 13158 4 _111_
rlabel metal2 s 9430 13056 9430 13056 4 _112_
rlabel metal1 s 10810 12852 10810 12852 4 _113_
rlabel metal2 s 11822 9724 11822 9724 4 _114_
rlabel metal1 s 11500 10234 11500 10234 4 _115_
rlabel metal1 s 12926 9690 12926 9690 4 _116_
rlabel metal1 s 12466 7752 12466 7752 4 _117_
rlabel metal2 s 13018 7990 13018 7990 4 _118_
rlabel metal2 s 14858 8194 14858 8194 4 _119_
rlabel metal1 s 14812 7786 14812 7786 4 _120_
rlabel metal2 s 15226 9588 15226 9588 4 _121_
rlabel metal1 s 13202 10013 13202 10013 4 _122_
rlabel metal1 s 13018 9554 13018 9554 4 _123_
rlabel metal1 s 13708 11186 13708 11186 4 _124_
rlabel metal2 s 13478 10506 13478 10506 4 _125_
rlabel metal1 s 12880 9146 12880 9146 4 _126_
rlabel metal2 s 14766 10931 14766 10931 4 _127_
rlabel metal2 s 14398 11730 14398 11730 4 _128_
rlabel metal1 s 14043 13158 14043 13158 4 _129_
rlabel metal2 s 13478 13090 13478 13090 4 _130_
rlabel metal1 s 15318 12818 15318 12818 4 _131_
rlabel metal1 s 14858 13226 14858 13226 4 _132_
rlabel metal1 s 16744 11594 16744 11594 4 _133_
rlabel metal1 s 16008 12818 16008 12818 4 _134_
rlabel metal1 s 16054 12886 16054 12886 4 _135_
rlabel metal2 s 14582 13770 14582 13770 4 _136_
rlabel metal1 s 13524 9894 13524 9894 4 _137_
rlabel metal2 s 15778 7616 15778 7616 4 _138_
rlabel metal1 s 11270 12886 11270 12886 4 _139_
rlabel metal1 s 8096 10030 8096 10030 4 _140_
rlabel metal1 s 6716 14042 6716 14042 4 _141_
rlabel metal1 s 4462 11152 4462 11152 4 _142_
rlabel metal1 s 7682 5338 7682 5338 4 _143_
rlabel metal1 s 9936 3366 9936 3366 4 _144_
rlabel metal2 s 13570 2992 13570 2992 4 _145_
rlabel metal1 s 12926 3706 12926 3706 4 _146_
rlabel metal2 s 9062 3910 9062 3910 4 _147_
rlabel metal2 s 6486 3264 6486 3264 4 _148_
rlabel metal2 s 1978 6154 1978 6154 4 _149_
rlabel metal1 s 10488 8602 10488 8602 4 _150_
rlabel metal2 s 9430 5134 9430 5134 4 _151_
rlabel metal1 s 2530 5712 2530 5712 4 _152_
rlabel metal2 s 3082 5916 3082 5916 4 _153_
rlabel metal1 s 9338 7820 9338 7820 4 _154_
rlabel metal1 s 7360 3706 7360 3706 4 _155_
rlabel metal1 s 9568 7854 9568 7854 4 _156_
rlabel metal2 s 12374 11424 12374 11424 4 _157_
rlabel metal1 s 11868 4250 11868 4250 4 _158_
rlabel metal1 s 10488 4250 10488 4250 4 _159_
rlabel metal2 s 10350 5236 10350 5236 4 _160_
rlabel metal1 s 8004 5270 8004 5270 4 _161_
rlabel metal1 s 10166 6800 10166 6800 4 _162_
rlabel metal2 s 9982 6868 9982 6868 4 _163_
rlabel metal2 s 10718 8738 10718 8738 4 _164_
rlabel metal1 s 9982 12750 9982 12750 4 _165_
rlabel metal1 s 13892 12070 13892 12070 4 _166_
rlabel metal2 s 15410 11594 15410 11594 4 _167_
rlabel metal2 s 3266 1027 3266 1027 4 clk
rlabel metal2 s 12466 9503 12466 9503 4 clknet_0_clk
rlabel metal1 s 8326 2890 8326 2890 4 clknet_2_0__leaf_clk
rlabel metal1 s 1840 7854 1840 7854 4 clknet_2_1__leaf_clk
rlabel metal1 s 14122 7412 14122 7412 4 clknet_2_2__leaf_clk
rlabel metal2 s 12926 14144 12926 14144 4 clknet_2_3__leaf_clk
rlabel metal3 s 0 10208 800 10328 4 count[0]
port 4 nsew
rlabel metal2 s 11638 1520 11638 1520 4 count[10]
rlabel metal2 s 10994 1520 10994 1520 4 count[11]
rlabel metal1 s 8510 3366 8510 3366 4 count[12]
rlabel metal2 s 10350 1520 10350 1520 4 count[13]
rlabel metal2 s 7774 1520 7774 1520 4 count[14]
rlabel metal2 s 9062 1520 9062 1520 4 count[15]
rlabel metal3 s 1096 12308 1096 12308 4 count[16]
rlabel metal3 s 0 11568 800 11688 4 count[17]
port 12 nsew
rlabel metal3 s 0 12928 800 13048 4 count[18]
port 13 nsew
rlabel metal3 s 0 14288 800 14408 4 count[19]
port 14 nsew
rlabel metal3 s 1372 8228 1372 8228 4 count[1]
rlabel metal2 s 9246 19839 9246 19839 4 count[20]
rlabel metal2 s 8602 19839 8602 19839 4 count[21]
rlabel metal1 s 11040 18938 11040 18938 4 count[22]
rlabel metal2 s 11914 19839 11914 19839 4 count[23]
rlabel metal2 s 17710 8857 17710 8857 4 count[24]
rlabel metal2 s 17710 8279 17710 8279 4 count[25]
rlabel metal2 s 17710 9503 17710 9503 4 count[26]
rlabel metal2 s 17710 10353 17710 10353 4 count[27]
rlabel metal2 s 17710 13855 17710 13855 4 count[28]
rlabel metal2 s 17710 14297 17710 14297 4 count[29]
rlabel metal3 s 0 7488 800 7608 4 count[2]
port 26 nsew
rlabel metal2 s 17710 13073 17710 13073 4 count[30]
rlabel metal3 s 17994 12308 17994 12308 4 count[31]
rlabel metal3 s 1326 6868 1326 6868 4 count[3]
rlabel metal2 s 5842 1520 5842 1520 4 count[4]
rlabel metal2 s 6486 1520 6486 1520 4 count[5]
rlabel metal2 s 7130 1520 7130 1520 4 count[6]
rlabel metal2 s 9706 1520 9706 1520 4 count[7]
rlabel metal2 s 12282 1656 12282 1656 4 count[8]
rlabel metal2 s 12926 1520 12926 1520 4 count[9]
rlabel metal3 s 1050 13668 1050 13668 4 en
rlabel metal2 s 2165 9554 2165 9554 4 net1
rlabel metal1 s 3634 12818 3634 12818 4 net10
rlabel metal1 s 1702 11764 1702 11764 4 net11
rlabel metal1 s 3174 13294 3174 13294 4 net12
rlabel metal2 s 4830 14212 4830 14212 4 net13
rlabel metal2 s 3174 8262 3174 8262 4 net14
rlabel metal1 s 9522 18734 9522 18734 4 net15
rlabel metal1 s 9108 13906 9108 13906 4 net16
rlabel metal2 s 8970 13736 8970 13736 4 net17
rlabel metal1 s 9522 11628 9522 11628 4 net18
rlabel metal1 s 14306 8432 14306 8432 4 net19
rlabel metal1 s 12650 4488 12650 4488 4 net2
rlabel metal1 s 17480 8466 17480 8466 4 net20
rlabel metal2 s 17526 9350 17526 9350 4 net21
rlabel metal2 s 17618 10438 17618 10438 4 net22
rlabel metal1 s 17043 13906 17043 13906 4 net23
rlabel metal1 s 15870 14042 15870 14042 4 net24
rlabel metal1 s 2208 5678 2208 5678 4 net25
rlabel metal2 s 17526 13022 17526 13022 4 net26
rlabel metal1 s 17480 11662 17480 11662 4 net27
rlabel metal1 s 2024 6766 2024 6766 4 net28
rlabel metal1 s 6164 2958 6164 2958 4 net29
rlabel metal1 s 1978 7820 1978 7820 4 net3
rlabel metal1 s 6394 2414 6394 2414 4 net30
rlabel metal1 s 7038 3366 7038 3366 4 net31
rlabel metal1 s 9292 2550 9292 2550 4 net32
rlabel metal1 s 12558 2414 12558 2414 4 net33
rlabel metal1 s 13938 4012 13938 4012 4 net34
rlabel metal1 s 1794 9622 1794 9622 4 net35
rlabel metal2 s 3634 7599 3634 7599 4 net36
rlabel metal1 s 12880 12206 12880 12206 4 net37
rlabel metal2 s 7590 7174 7590 7174 4 net38
rlabel metal1 s 8418 8874 8418 8874 4 net39
rlabel metal1 s 11960 2414 11960 2414 4 net4
rlabel metal1 s 11454 8840 11454 8840 4 net40
rlabel metal2 s 10350 9996 10350 9996 4 net41
rlabel metal1 s 6670 13362 6670 13362 4 net42
rlabel metal1 s 13340 13498 13340 13498 4 net43
rlabel metal1 s 15042 13328 15042 13328 4 net44
rlabel metal2 s 1518 7888 1518 7888 4 net45
rlabel metal1 s 9752 13770 9752 13770 4 net46
rlabel metal1 s 1656 9554 1656 9554 4 net47
rlabel metal1 s 8740 5338 8740 5338 4 net48
rlabel metal2 s 10258 3706 10258 3706 4 net49
rlabel metal1 s 10856 3162 10856 3162 4 net5
rlabel metal2 s 9154 3332 9154 3332 4 net50
rlabel metal1 s 16330 7378 16330 7378 4 net51
rlabel metal2 s 6762 14076 6762 14076 4 net52
rlabel metal1 s 13478 2448 13478 2448 4 net53
rlabel metal1 s 6578 3060 6578 3060 4 net54
rlabel metal1 s 15272 14382 15272 14382 4 net55
rlabel metal2 s 7314 5406 7314 5406 4 net56
rlabel metal1 s 13478 3502 13478 3502 4 net57
rlabel metal1 s 2300 9622 2300 9622 4 net58
rlabel metal1 s 8372 12750 8372 12750 4 net59
rlabel metal2 s 7958 4386 7958 4386 4 net6
rlabel metal1 s 9752 6290 9752 6290 4 net60
rlabel metal1 s 2484 6766 2484 6766 4 net61
rlabel metal1 s 16652 12818 16652 12818 4 net62
rlabel metal1 s 1748 7378 1748 7378 4 net63
rlabel metal1 s 3910 5236 3910 5236 4 net64
rlabel metal2 s 11730 12988 11730 12988 4 net65
rlabel metal1 s 4554 4080 4554 4080 4 net66
rlabel metal1 s 6026 10030 6026 10030 4 net67
rlabel metal1 s 10074 5542 10074 5542 4 net7
rlabel metal1 s 7820 2346 7820 2346 4 net8
rlabel metal1 s 8970 2414 8970 2414 4 net9
rlabel metal2 s 17802 4369 17802 4369 4 rst_n
flabel metal4 s 4868 2128 5188 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4208 2128 4528 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 3238 0 3294 800 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal3 s 400 10268 400 10268 0 FreeSans 600 0 0 0 count[0]
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 count[10]
port 5 nsew
flabel metal2 s 10966 0 11022 800 0 FreeSans 280 90 0 0 count[11]
port 6 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 count[12]
port 7 nsew
flabel metal2 s 10322 0 10378 800 0 FreeSans 280 90 0 0 count[13]
port 8 nsew
flabel metal2 s 7746 0 7802 800 0 FreeSans 280 90 0 0 count[14]
port 9 nsew
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 count[15]
port 10 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 count[16]
port 11 nsew
flabel metal3 s 400 11628 400 11628 0 FreeSans 600 0 0 0 count[17]
flabel metal3 s 400 12988 400 12988 0 FreeSans 600 0 0 0 count[18]
flabel metal3 s 400 14348 400 14348 0 FreeSans 600 0 0 0 count[19]
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 count[1]
port 15 nsew
flabel metal2 s 9034 20648 9090 21448 0 FreeSans 280 90 0 0 count[20]
port 16 nsew
flabel metal2 s 8390 20648 8446 21448 0 FreeSans 280 90 0 0 count[21]
port 17 nsew
flabel metal2 s 10966 20648 11022 21448 0 FreeSans 280 90 0 0 count[22]
port 18 nsew
flabel metal2 s 11610 20648 11666 21448 0 FreeSans 280 90 0 0 count[23]
port 19 nsew
flabel metal3 s 18504 8848 19304 8968 0 FreeSans 600 0 0 0 count[24]
port 20 nsew
flabel metal3 s 18504 8168 19304 8288 0 FreeSans 600 0 0 0 count[25]
port 21 nsew
flabel metal3 s 18504 9528 19304 9648 0 FreeSans 600 0 0 0 count[26]
port 22 nsew
flabel metal3 s 18504 10208 19304 10328 0 FreeSans 600 0 0 0 count[27]
port 23 nsew
flabel metal3 s 18504 13608 19304 13728 0 FreeSans 600 0 0 0 count[28]
port 24 nsew
flabel metal3 s 18504 14288 19304 14408 0 FreeSans 600 0 0 0 count[29]
port 25 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 count[2]
flabel metal3 s 18504 12928 19304 13048 0 FreeSans 600 0 0 0 count[30]
port 27 nsew
flabel metal3 s 18504 12248 19304 12368 0 FreeSans 600 0 0 0 count[31]
port 28 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 count[3]
port 29 nsew
flabel metal2 s 5814 0 5870 800 0 FreeSans 280 90 0 0 count[4]
port 30 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 count[5]
port 31 nsew
flabel metal2 s 7102 0 7158 800 0 FreeSans 280 90 0 0 count[6]
port 32 nsew
flabel metal2 s 9678 0 9734 800 0 FreeSans 280 90 0 0 count[7]
port 33 nsew
flabel metal2 s 12254 0 12310 800 0 FreeSans 280 90 0 0 count[8]
port 34 nsew
flabel metal2 s 12898 0 12954 800 0 FreeSans 280 90 0 0 count[9]
port 35 nsew
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 en
port 36 nsew
flabel metal3 s 18504 4088 19304 4208 0 FreeSans 600 0 0 0 rst_n
port 37 nsew
<< properties >>
string FIXED_BBOX 0 0 140000 140000
<< end >>
