* NGSPICE file created from counter32.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

.subckt counter32 VGND VPWR clk count[0] count[10] count[11] count[12] count[13] count[14]
+ count[15] count[16] count[17] count[18] count[19] count[1] count[20] count[21] count[22]
+ count[23] count[24] count[25] count[26] count[27] count[28] count[29] count[2] count[30]
+ count[31] count[3] count[4] count[5] count[6] count[7] count[8] count[9] en rst_n
XTAP_TAPCELL_ROW_24_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_294_ _045_ _094_ _124_ net43 VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__o31ai_1
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_363_ clknet_2_3__leaf_clk _027_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfxtp_1
XFILLER_3_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_346_ clknet_2_2__leaf_clk _010_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfxtp_1
X_277_ _165_ _054_ _112_ _039_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__nand4_1
X_200_ _055_ _057_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_4_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_329_ net31 net30 VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__and2_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput20 net20 VGND VGND VPWR VPWR count[25] sky130_fd_sc_hd__buf_2
Xoutput7 net7 VGND VGND VPWR VPWR count[13] sky130_fd_sc_hd__buf_2
Xoutput31 net31 VGND VGND VPWR VPWR count[6] sky130_fd_sc_hd__buf_2
XFILLER_22_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_293_ net27 net26 _166_ _035_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__a31o_1
X_362_ clknet_2_3__leaf_clk _026_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfxtp_1
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_276_ net17 net16 net15 net46 VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_20_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_345_ clknet_2_2__leaf_clk _009_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259_ _046_ net39 net41 _038_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__nand4_1
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_328_ net28 net25 net14 net3 VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__nand4_4
XFILLER_15_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold20 net11 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 net10 VGND VGND VPWR VPWR count[16] sky130_fd_sc_hd__buf_2
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput21 net21 VGND VGND VPWR VPWR count[26] sky130_fd_sc_hd__buf_2
Xoutput32 net32 VGND VGND VPWR VPWR count[7] sky130_fd_sc_hd__buf_2
Xoutput8 net8 VGND VGND VPWR VPWR count[14] sky130_fd_sc_hd__buf_2
XFILLER_22_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_292_ _121_ _123_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nor2_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_361_ clknet_2_2__leaf_clk _025_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfxtp_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_275_ _043_ _094_ net17 VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_11_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ clknet_2_2__leaf_clk _008_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_189_ net17 net16 net15 VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__and3_1
X_258_ _050_ net39 net10 net41 net67 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__a41oi_1
X_327_ net28 net25 _152_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__and3_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold10 net34 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput11 net11 VGND VGND VPWR VPWR count[17] sky130_fd_sc_hd__buf_2
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput22 net22 VGND VGND VPWR VPWR count[27] sky130_fd_sc_hd__buf_2
XFILLER_15_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput33 net33 VGND VGND VPWR VPWR count[8] sky130_fd_sc_hd__buf_2
Xoutput9 net9 VGND VGND VPWR VPWR count[15] sky130_fd_sc_hd__buf_2
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_291_ _034_ _114_ net43 VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__o21ai_1
X_360_ clknet_2_2__leaf_clk _024_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfxtp_2
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_274_ _110_ _109_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__nor2_1
X_343_ clknet_2_0__leaf_clk _007_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfxtp_1
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_188_ _036_ _039_ _041_ _044_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__nand4_2
X_257_ _097_ _098_ net42 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__and3_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_326_ net14 net3 VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_8_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_309_ net62 VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__inv_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold11 net3 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_20_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput23 net23 VGND VGND VPWR VPWR count[28] sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR count[18] sky130_fd_sc_hd__buf_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput34 net34 VGND VGND VPWR VPWR count[9] sky130_fd_sc_hd__buf_2
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_290_ net40 _033_ _053_ _116_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__nand4_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_273_ _043_ _095_ net42 VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__o21ai_1
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_342_ clknet_2_0__leaf_clk _006_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_187_ _039_ _041_ _044_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__nand3_1
X_256_ _046_ net39 net10 net41 VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__nand4_1
X_325_ net42 VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__inv_2
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
X_308_ net27 _133_ net44 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__o21a_1
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_239_ _051_ net38 net6 VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__and3_1
XFILLER_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold12 net16 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR count[29] sky130_fd_sc_hd__buf_2
Xoutput13 net13 VGND VGND VPWR VPWR count[19] sky130_fd_sc_hd__buf_2
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_272_ _165_ _054_ _042_ net47 net59 VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__a41oi_1
XTAP_TAPCELL_ROW_20_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_341_ clknet_2_0__leaf_clk _005_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfxtp_1
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_186_ net18 net17 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__and2_1
XFILLER_13_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_255_ _050_ net39 net41 net10 VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__a31o_1
X_324_ net46 VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__inv_2
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_2
X_307_ _135_ _131_ _134_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__a21oi_1
X_169_ net9 net8 net7 net6 VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__nand4_2
X_238_ _051_ net38 net6 VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold13 net7 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput25 net25 VGND VGND VPWR VPWR count[2] sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR count[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_23_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_271_ _140_ _105_ net42 _108_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__o211a_1
XFILLER_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_340_ clknet_2_0__leaf_clk _004_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_185_ _039_ _041_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__nand2_1
X_254_ _143_ _092_ _096_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a21oi_1
X_323_ net61 VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_306_ _167_ _127_ _128_ net44 VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__o31ai_1
X_237_ _144_ _080_ _083_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__a21oi_1
X_168_ net7 net6 VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__nand2_1
XFILLER_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold14 net28 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput15 net15 VGND VGND VPWR VPWR count[20] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput26 net26 VGND VGND VPWR VPWR count[30] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_270_ _140_ _106_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__nand2_1
XFILLER_5_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_322_ net54 VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__inv_2
X_184_ net15 net13 net12 _038_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and4_1
X_253_ _050_ net39 net41 _151_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_305_ _167_ _127_ _128_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__nor3_1
X_236_ net36 _082_ _151_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__a21o_1
XFILLER_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold15 net26 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_219_ _070_ net42 VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput16 net16 VGND VGND VPWR VPWR count[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput27 net27 VGND VGND VPWR VPWR count[31] sky130_fd_sc_hd__buf_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_183_ net16 net15 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__and2_1
X_252_ _050_ net39 net41 VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__nand3_1
X_321_ net50 VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_304_ _136_ _130_ _132_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_3_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_235_ _150_ _154_ _156_ _160_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nor4_1
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold16 net14 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_218_ net35 _065_ net45 _155_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_6_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput17 net17 VGND VGND VPWR VPWR count[22] sky130_fd_sc_hd__buf_2
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput28 net28 VGND VGND VPWR VPWR count[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_182_ net13 net12 net11 net10 VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand4_2
X_251_ net46 _157_ _164_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__nand3_1
Xfanout41 _164_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_320_ net57 VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__inv_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_303_ _131_ net44 VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__nand2_1
X_234_ _145_ _078_ _081_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold17 net29 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_217_ _067_ _069_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__nor2_1
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput18 net18 VGND VGND VPWR VPWR count[23] sky130_fd_sc_hd__buf_2
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput29 net29 VGND VGND VPWR VPWR count[4] sky130_fd_sc_hd__buf_2
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_181_ net13 net12 net11 net10 VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__and4_2
Xfanout42 net44 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
X_250_ _091_ _093_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ net40 _166_ _053_ net37 VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__nand4_1
X_233_ _080_ net43 VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__nand2_1
Xhold18 net18 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_216_ _068_ net42 VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__nand2_1
XFILLER_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput19 net19 VGND VGND VPWR VPWR count[24] sky130_fd_sc_hd__buf_2
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_180_ net11 net10 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__and2_1
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout43 net44 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_301_ _130_ net43 _129_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and3_1
X_232_ net36 _159_ _157_ net46 VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__nand4_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold19 net30 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_7_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_215_ net35 _065_ net30 net45 VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__nand4_1
XFILLER_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap40 _165_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout44 net2 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_300_ net23 net40 _049_ net37 VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__nand4_1
X_231_ _146_ _076_ _079_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_23_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput1 en VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_214_ net35 _065_ net45 net66 VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__a31oi_1
XFILLER_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout45 net47 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
XFILLER_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_230_ _078_ net43 VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__nand2_1
X_359_ clknet_2_3__leaf_clk _023_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfxtp_1
Xinput2 rst_n VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_213_ _064_ _066_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__nor2_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout46 net47 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xfanout35 net36 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
XFILLER_5_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_358_ clknet_2_3__leaf_clk _022_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ _056_ _119_ net21 VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__o21ba_1
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_212_ net35 _065_ net45 _151_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__a31o_1
XFILLER_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout47 net1 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
Xfanout36 _051_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_357_ clknet_2_1__leaf_clk _021_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_1_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_288_ _138_ _118_ _120_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_211_ net29 net28 net25 _152_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_27_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_356_ clknet_2_3__leaf_clk _020_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfxtp_1
X_287_ _056_ _119_ net43 VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_210_ net35 _153_ net45 net64 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__a31oi_1
X_339_ clknet_2_0__leaf_clk _003_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_355_ clknet_2_1__leaf_clk _019_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfxtp_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_286_ _032_ _035_ net20 net19 net46 VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__o2111ai_2
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_269_ _141_ _104_ _107_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a21oi_1
X_338_ clknet_2_1__leaf_clk _002_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfxtp_1
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_354_ clknet_2_1__leaf_clk _018_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_1
X_285_ _117_ _118_ net43 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__and3_1
XFILLER_30_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_268_ _040_ _095_ net42 VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__o21ai_1
X_199_ net35 net47 net3 _151_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__a31o_1
XFILLER_2_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_337_ clknet_2_1__leaf_clk _001_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfxtp_1
XFILLER_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_284_ net19 net40 _053_ _116_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__nand4_1
XFILLER_14_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_353_ clknet_2_1__leaf_clk _017_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_198_ _157_ _164_ _047_ _052_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__nand4_2
X_267_ _050_ net39 net41 _039_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__nand4_1
X_336_ clknet_2_1__leaf_clk _000_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfxtp_2
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_319_ net53 VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__inv_2
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_352_ clknet_2_1__leaf_clk _016_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_2
X_283_ _150_ _056_ net19 VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__o21bai_1
XFILLER_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_266_ _046_ net39 net41 _039_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__nand4_1
X_197_ net35 net47 net58 VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__a21oi_1
X_335_ net7 net6 VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_22_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap38 _082_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_318_ net49 VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__inv_2
X_249_ _092_ net42 VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_30_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 net9 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_282_ _139_ _113_ _115_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__a21oi_1
X_351_ clknet_2_0__leaf_clk _015_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfxtp_1
XFILLER_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_334_ net5 net4 net34 net33 VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_19_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_196_ net18 _036_ _039_ _047_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__nand4_1
X_265_ _142_ _100_ net42 _102_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__o211a_1
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap39 _072_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_16_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_248_ net36 net38 net8 _161_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_317_ net48 VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__inv_2
X_179_ _032_ _035_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__or2_1
XFILLER_20_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2 net5 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_281_ _137_ _032_ _034_ net47 VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__o31a_1
X_350_ clknet_2_0__leaf_clk _014_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfxtp_1
XFILLER_19_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_264_ net47 _165_ _054_ _103_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__nand4_1
X_195_ _139_ _040_ _047_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__nor3b_1
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ net4 net34 net33 VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__and3_1
X_316_ net12 VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_247_ _051_ net38 _161_ net56 VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_7_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_178_ _032_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nor2_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 net32 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_280_ _114_ net43 VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__nand2_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_263_ net12 net11 net10 VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__and3_1
X_194_ _139_ _040_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__nor2_1
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_332_ net34 net33 VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_26_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_315_ net52 VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__inv_2
X_177_ net22 net21 net20 net19 VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nand4_4
X_246_ _086_ _090_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_21_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ net36 _158_ _157_ net46 VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__nand4_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 net20 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_29_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_262_ _142_ _101_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__nand2_1
X_193_ _157_ _164_ _036_ _049_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__nand4_2
X_331_ _154_ _156_ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__nor2_4
XFILLER_17_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_176_ net21 net20 net19 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nand3_1
X_314_ net15 VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__inv_2
X_245_ _089_ net43 VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__nand2_1
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_228_ _074_ _077_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__nor2_1
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 net13 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_192_ _036_ _049_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__nand2_2
X_261_ _151_ _099_ _100_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__nor3b_1
X_330_ net32 net31 net30 net29 VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__nand4_4
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_313_ net65 VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__inv_2
X_175_ net21 net20 net19 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__and3_1
X_244_ _037_ _056_ _088_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__o21bai_1
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ _076_ net43 VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__nand2_1
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 net4 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_260_ _050_ net39 net41 _038_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__nand4_1
X_191_ _040_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nor2_2
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_174_ net27 net26 net24 net23 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nand4_4
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_243_ net46 _157_ _087_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__nand3_1
X_312_ net51 VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_226_ _037_ _056_ _075_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 net31 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_209_ _149_ _061_ _063_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_190_ net18 net17 net16 net15 VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__nand4_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_173_ net26 _166_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__nand2_1
X_311_ net22 VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__inv_2
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_242_ _160_ _162_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__nor2_1
XFILLER_11_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_225_ net33 net46 _157_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 net24 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
X_208_ net35 _153_ net45 _151_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_5_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_310_ net55 VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__inv_2
XFILLER_11_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_172_ net24 net23 VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_15_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_241_ net36 _082_ net6 net60 VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_30_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_224_ net36 _157_ net46 net33 VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__a31oi_1
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 net8 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_207_ _060_ _062_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_171_ _154_ _156_ _160_ _163_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__nor4_2
X_240_ _151_ _084_ _085_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_30_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_223_ _147_ _070_ _073_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_206_ _061_ net42 VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nand2_1
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_170_ _160_ _163_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_30_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_299_ _127_ _128_ net23 VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_15_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_222_ net36 _157_ net46 _151_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__a31o_1
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_205_ net35 _152_ net45 net25 VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__nand4_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_367_ clknet_2_3__leaf_clk _031_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
X_298_ _137_ _122_ _125_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_25_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_221_ _150_ _154_ _156_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nor3_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_204_ net36 _152_ net45 net25 VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__a31oi_1
XFILLER_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput3 net3 VGND VGND VPWR VPWR count[0] sky130_fd_sc_hd__buf_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_366_ clknet_2_3__leaf_clk _030_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfxtp_1
X_297_ _157_ _164_ _049_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__nand3_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire37 _126_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_12_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_220_ _148_ _068_ _071_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_0_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_349_ clknet_2_2__leaf_clk _013_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_203_ _058_ _059_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__nor2_1
XFILLER_9_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput4 net4 VGND VGND VPWR VPWR count[10] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_365_ clknet_2_3__leaf_clk _029_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfxtp_1
X_296_ _032_ _033_ net22 net47 VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__nand4_1
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_279_ _032_ _035_ _049_ _072_ net41 VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__o2111ai_2
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_348_ clknet_2_1__leaf_clk _012_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfxtp_1
XFILLER_17_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_202_ net36 _152_ net45 _151_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__a31o_1
XFILLER_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput5 net5 VGND VGND VPWR VPWR count[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_364_ clknet_2_3__leaf_clk _028_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfxtp_1
X_295_ _137_ _150_ _034_ _032_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__nor4b_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_278_ _113_ net44 _111_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__and3_1
X_347_ clknet_2_0__leaf_clk _011_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfxtp_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_201_ net35 net45 net3 net63 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__a31oi_1
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput6 net6 VGND VGND VPWR VPWR count[12] sky130_fd_sc_hd__buf_2
Xoutput30 net30 VGND VGND VPWR VPWR count[5] sky130_fd_sc_hd__buf_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

